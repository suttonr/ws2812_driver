// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Fri Nov 28 22:57:04 2025
//
// Verilog Description of module top
//

module top (sclk, sclk_enable, ws2813_out, MISO_SLAVE, MOSI_SLAVE, 
            CSn_SLAVE, SCLK_SLAVE, SPI_RST, led0, led1, led2, led3, 
            led4, led5, led6, led7, yled0, yled1, yled2, yled3, 
            yled4, yled5, yled6, yled7);   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(6[8:11])
    input sclk;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    output sclk_enable;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(9[3:14])
    output [20:0]ws2813_out;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    output MISO_SLAVE;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(13[6:16])
    input MOSI_SLAVE;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(14[9:19])
    input CSn_SLAVE;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(15[9:18])
    input SCLK_SLAVE;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(16[9:19])
    input SPI_RST;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(17[3:10])
    output led0 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[3:7])
    output led1 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[8:12])
    output led2 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[13:17])
    output led3 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[18:22])
    output led4 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[23:27])
    output led5 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[28:32])
    output led6 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[33:37])
    input led7 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[38:42])
    output yled0 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[3:8])
    output yled1 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[9:14])
    output yled2 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[15:20])
    output yled3 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[21:26])
    output yled4 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[27:32])
    output yled5 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[33:38])
    output yled6 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[39:44])
    input yled7 /* synthesis .original_dir=IN_OUT */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[45:50])
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire SCLK_SLAVE_c /* synthesis is_clock=1, SET_AS_NETWORK=SCLK_SLAVE_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(16[9:19])
    
    wire GND_net, VCC_net, ws2813_out_c_20, ws2813_out_c_19, ws2813_out_c_18, 
        ws2813_out_c_17, ws2813_out_c_16, ws2813_out_c_15, ws2813_out_c_14, 
        ws2813_out_c_13, ws2813_out_c_12, ws2813_out_c_11, ws2813_out_c_10, 
        ws2813_out_c_9, ws2813_out_c_8, ws2813_out_c_7, ws2813_out_c_6, 
        ws2813_out_c_5, ws2813_out_c_4, ws2813_out_c_3, ws2813_out_c_2, 
        ws2813_out_c_1, ws2813_out_c_0, MOSI_SLAVE_c, CSn_SLAVE_c, SPI_RST_c, 
        yled0_c, yled1_c, yled2_c, yled3_c, yled4_c, yled5_c, yled6_c;
    wire [8:0]WrAddress;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(96[12:21])
    wire [8:0]\RdAddress[0] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[1] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[2] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[3] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[4] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[5] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[6] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[7] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[8] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[9] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[10] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[11] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[12] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[13] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[14] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[15] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[16] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[17] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[18] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[19] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [8:0]\RdAddress[20] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(97[9:18])
    wire [23:0]Data;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(98[12:16])
    wire [23:0]WE;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(99[12:14])
    wire [23:0]\Q[0] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[1] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[2] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[3] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[4] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[5] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[6] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[7] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[8] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[9] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[10] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[11] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[12] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[13] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[14] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[15] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[16] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[17] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[18] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[19] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [23:0]\Q[20] ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(103[9:10])
    wire [0:20]port_status;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(104[9:20])
    
    wire CSn;
    wire [7:0]DATA_OUT;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(111[12:20])
    
    wire RX_RDY;
    wire [5:0]rx_data_cnt;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(91[25:36])
    
    wire rx_data_cnt_5__N_63;
    wire [2:0]state_adj_1050;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    wire [2:0]state_adj_1482;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    wire [2:0]state_adj_1590;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire n13101, n10470, n41629, n54591, n54583, n34568, SCLK_SLAVE_c_enable_5, 
        n50005;
    
    VHI i2 (.Z(VCC_net));
    \WS2812(48000000,"111111111")  WS2812_9 (.sclk_c(sclk_c), .\port_status[9] (port_status[9]), 
            .ws2813_out_c_9(ws2813_out_c_9), .GND_net(GND_net), .\Q[9] ({\Q[9] }), 
            .\RdAddress[9] ({\RdAddress[9] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(234[12:18])
    frame_buffer_0_U9 framebuffer19 (.WrAddress({WrAddress}), .\RdAddress[19] ({\RdAddress[19] }), 
            .Data({Data}), .\WE[19] (WE[19]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[19] ({\Q[19] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(339[17:31])
    frame_buffer_0_U7 framebuffer20 (.WrAddress({WrAddress}), .\RdAddress[20] ({\RdAddress[20] }), 
            .Data({Data}), .\WE[20] (WE[20]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[20] ({\Q[20] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(350[17:31])
    frame_buffer_0_U6 framebuffer2 (.WrAddress({WrAddress}), .\RdAddress[2] ({\RdAddress[2] }), 
            .Data({Data}), .\WE[2] (WE[2]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[2] ({\Q[2] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(152[16:30])
    frame_buffer_0_U5 framebuffer3 (.WrAddress({WrAddress}), .\RdAddress[3] ({\RdAddress[3] }), 
            .Data({Data}), .\WE[3] (WE[3]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[3] ({\Q[3] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(163[16:30])
    frame_buffer_0_U4 framebuffer4 (.WrAddress({WrAddress}), .\RdAddress[4] ({\RdAddress[4] }), 
            .Data({Data}), .\WE[4] (WE[4]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[4] ({\Q[4] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(174[16:30])
    frame_buffer_0_U3 framebuffer5 (.WrAddress({WrAddress}), .\RdAddress[5] ({\RdAddress[5] }), 
            .Data({Data}), .\WE[5] (WE[5]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[5] ({\Q[5] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(185[16:30])
    frame_buffer_0_U2 framebuffer6 (.WrAddress({WrAddress}), .\RdAddress[6] ({\RdAddress[6] }), 
            .Data({Data}), .\WE[6] (WE[6]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[6] ({\Q[6] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(196[16:30])
    frame_buffer_0_U1 framebuffer7 (.WrAddress({WrAddress}), .\RdAddress[7] ({\RdAddress[7] }), 
            .Data({Data}), .\WE[7] (WE[7]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[7] ({\Q[7] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(207[16:30])
    frame_buffer_0_U0 framebuffer8 (.WrAddress({WrAddress}), .\RdAddress[8] ({\RdAddress[8] }), 
            .Data({Data}), .\WE[8] (WE[8]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[8] ({\Q[8] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(218[16:30])
    frame_buffer_0_U19 framebuffer0 (.WrAddress({WrAddress}), .\RdAddress[0] ({\RdAddress[0] }), 
            .Data({Data}), .\WE[0] (WE[0]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[0] ({\Q[0] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(130[16:30])
    frame_buffer_0_U18 framebuffer10 (.WrAddress({WrAddress}), .\RdAddress[10] ({\RdAddress[10] }), 
            .Data({Data}), .\WE[10] (WE[10]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[10] ({\Q[10] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(240[17:31])
    frame_buffer_0_U17 framebuffer11 (.WrAddress({WrAddress}), .\RdAddress[11] ({\RdAddress[11] }), 
            .Data({Data}), .\WE[11] (WE[11]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[11] ({\Q[11] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(251[17:31])
    frame_buffer_0_U16 framebuffer12 (.WrAddress({WrAddress}), .\RdAddress[12] ({\RdAddress[12] }), 
            .Data({Data}), .\WE[12] (WE[12]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[12] ({\Q[12] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(262[17:31])
    frame_buffer_0_U15 framebuffer13 (.WrAddress({WrAddress}), .\RdAddress[13] ({\RdAddress[13] }), 
            .Data({Data}), .\WE[13] (WE[13]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[13] ({\Q[13] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(273[17:31])
    frame_buffer_0_U14 framebuffer14 (.WrAddress({WrAddress}), .\RdAddress[14] ({\RdAddress[14] }), 
            .Data({Data}), .\WE[14] (WE[14]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[14] ({\Q[14] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(284[17:31])
    frame_buffer_0_U13 framebuffer15 (.WrAddress({WrAddress}), .\RdAddress[15] ({\RdAddress[15] }), 
            .Data({Data}), .\WE[15] (WE[15]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[15] ({\Q[15] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(295[17:31])
    frame_buffer_0_U12 framebuffer16 (.WrAddress({WrAddress}), .\RdAddress[16] ({\RdAddress[16] }), 
            .Data({Data}), .\WE[16] (WE[16]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[16] ({\Q[16] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(306[17:31])
    frame_buffer_0_U11 framebuffer17 (.WrAddress({WrAddress}), .\RdAddress[17] ({\RdAddress[17] }), 
            .Data({Data}), .\WE[17] (WE[17]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[17] ({\Q[17] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(317[17:31])
    frame_buffer_0_U10 framebuffer18 (.WrAddress({WrAddress}), .\RdAddress[18] ({\RdAddress[18] }), 
            .Data({Data}), .\WE[18] (WE[18]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[18] ({\Q[18] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(328[17:31])
    frame_buffer_0_U8 framebuffer1 (.WrAddress({WrAddress}), .\RdAddress[1] ({\RdAddress[1] }), 
            .Data({Data}), .\WE[1] (WE[1]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[1] ({\Q[1] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(141[16:30])
    OB sclk_enable_pad (.I(VCC_net), .O(sclk_enable));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(9[3:14])
    LUT4 i29232_2_lut_rep_580_3_lut (.A(state_adj_1590[0]), .B(state_adj_1590[2]), 
         .C(state_adj_1590[1]), .Z(n54583)) /* synthesis lut_function=(A+(B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(18[3:9])
    defparam i29232_2_lut_rep_580_3_lut.init = 16'heaea;
    LUT4 i29947_2_lut_rep_588_3_lut (.A(state_adj_1482[0]), .B(state_adj_1482[2]), 
         .C(state_adj_1482[1]), .Z(n54591)) /* synthesis lut_function=(A+(B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(18[3:9])
    defparam i29947_2_lut_rep_588_3_lut.init = 16'heaea;
    OB ws2813_out_pad_20 (.I(ws2813_out_c_20), .O(ws2813_out[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_19 (.I(ws2813_out_c_19), .O(ws2813_out[19]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_18 (.I(ws2813_out_c_18), .O(ws2813_out[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_17 (.I(ws2813_out_c_17), .O(ws2813_out[17]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_16 (.I(ws2813_out_c_16), .O(ws2813_out[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_15 (.I(ws2813_out_c_15), .O(ws2813_out[15]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_14 (.I(ws2813_out_c_14), .O(ws2813_out[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_13 (.I(ws2813_out_c_13), .O(ws2813_out[13]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_12 (.I(ws2813_out_c_12), .O(ws2813_out[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_11 (.I(ws2813_out_c_11), .O(ws2813_out[11]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_10 (.I(ws2813_out_c_10), .O(ws2813_out[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_9 (.I(ws2813_out_c_9), .O(ws2813_out[9]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_8 (.I(ws2813_out_c_8), .O(ws2813_out[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_7 (.I(ws2813_out_c_7), .O(ws2813_out[7]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_6 (.I(ws2813_out_c_6), .O(ws2813_out[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_5 (.I(ws2813_out_c_5), .O(ws2813_out[5]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_4 (.I(ws2813_out_c_4), .O(ws2813_out[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_3 (.I(ws2813_out_c_3), .O(ws2813_out[3]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_2 (.I(ws2813_out_c_2), .O(ws2813_out[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_1 (.I(ws2813_out_c_1), .O(ws2813_out[1]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OB ws2813_out_pad_0 (.I(ws2813_out_c_0), .O(ws2813_out[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(10[3:13])
    OBZ MISO_SLAVE_pad (.I(GND_net), .T(CSn_SLAVE_c), .O(MISO_SLAVE));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(341[14] 351[26])
    OB led0_pad (.I(VCC_net), .O(led0));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[3:7])
    OB led1_pad (.I(VCC_net), .O(led1));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[8:12])
    OB led2_pad (.I(VCC_net), .O(led2));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[13:17])
    OB led3_pad (.I(VCC_net), .O(led3));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[18:22])
    OB led4_pad (.I(VCC_net), .O(led4));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[23:27])
    OB led5_pad (.I(VCC_net), .O(led5));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[28:32])
    OB led6_pad (.I(VCC_net), .O(led6));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(21[33:37])
    OB yled0_pad (.I(yled0_c), .O(yled0));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[3:8])
    OB yled1_pad (.I(yled1_c), .O(yled1));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[9:14])
    OB yled2_pad (.I(yled2_c), .O(yled2));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[15:20])
    OB yled3_pad (.I(yled3_c), .O(yled3));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[21:26])
    OB yled4_pad (.I(yled4_c), .O(yled4));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[27:32])
    OB yled5_pad (.I(yled5_c), .O(yled5));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[33:38])
    OB yled6_pad (.I(yled6_c), .O(yled6));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(23[39:44])
    IB sclk_pad (.I(sclk), .O(sclk_c));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    IB MOSI_SLAVE_pad (.I(MOSI_SLAVE), .O(MOSI_SLAVE_c));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(14[9:19])
    IB CSn_SLAVE_pad (.I(CSn_SLAVE), .O(CSn_SLAVE_c));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(15[9:18])
    IB SCLK_SLAVE_pad (.I(SCLK_SLAVE), .O(SCLK_SLAVE_c));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(16[9:19])
    IB SPI_RST_pad (.I(SPI_RST), .O(SPI_RST_c));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(17[3:10])
    LUT4 i29460_2_lut_3_lut (.A(state_adj_1050[0]), .B(state_adj_1050[2]), 
         .C(state_adj_1050[1]), .Z(n41629)) /* synthesis lut_function=(A+(B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(18[3:9])
    defparam i29460_2_lut_3_lut.init = 16'heaea;
    LUT4 i38441_2_lut_rep_679 (.A(CSn_SLAVE_c), .B(rx_data_cnt_5__N_63), 
         .Z(SCLK_SLAVE_c_enable_5)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i38441_2_lut_rep_679.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut (.A(CSn_SLAVE_c), .B(rx_data_cnt_5__N_63), .C(rx_data_cnt[0]), 
         .Z(n50005)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2d2d;
    LUT4 state_2__bdd_4_lut (.A(state_adj_1050[2]), .B(state_adj_1050[0]), 
         .C(n13101), .D(state_adj_1050[1]), .Z(n10470)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (C (D))) */ ;
    defparam state_2__bdd_4_lut.init = 16'hfa80;
    LUT4 i22356_1_lut (.A(SPI_RST_c), .Z(n34568)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(17[3:10])
    defparam i22356_1_lut.init = 16'h5555;
    LUT4 i2_3_lut (.A(port_status[2]), .B(port_status[1]), .C(port_status[0]), 
         .Z(yled0_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(383[11:61])
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_adj_928 (.A(port_status[5]), .B(port_status[4]), .C(port_status[3]), 
         .Z(yled1_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(384[14:64])
    defparam i2_3_lut_adj_928.init = 16'hfefe;
    LUT4 i2_3_lut_adj_929 (.A(port_status[8]), .B(port_status[7]), .C(port_status[6]), 
         .Z(yled2_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(385[14:64])
    defparam i2_3_lut_adj_929.init = 16'hfefe;
    LUT4 i2_3_lut_adj_930 (.A(port_status[11]), .B(port_status[10]), .C(port_status[9]), 
         .Z(yled3_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(386[14:66])
    defparam i2_3_lut_adj_930.init = 16'hfefe;
    LUT4 i2_3_lut_adj_931 (.A(port_status[14]), .B(port_status[13]), .C(port_status[12]), 
         .Z(yled4_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(387[14:67])
    defparam i2_3_lut_adj_931.init = 16'hfefe;
    LUT4 i2_3_lut_adj_932 (.A(port_status[17]), .B(port_status[16]), .C(port_status[15]), 
         .Z(yled5_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(388[14:67])
    defparam i2_3_lut_adj_932.init = 16'hfefe;
    LUT4 i2_3_lut_adj_933 (.A(port_status[20]), .B(port_status[19]), .C(port_status[18]), 
         .Z(yled6_c)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(389[14:67])
    defparam i2_3_lut_adj_933.init = 16'hfefe;
    \load_mem(48000000)  load_mem_t (.GND_net(GND_net), .Data({Data}), .sclk_c(sclk_c), 
            .CSn(CSn), .WrAddress({WrAddress}), .\WE[0] (WE[0]), .DATA_OUT({DATA_OUT}), 
            .RX_RDY(RX_RDY), .\WE[1] (WE[1]), .\WE[2] (WE[2]), .\WE[3] (WE[3]), 
            .\WE[4] (WE[4]), .\WE[5] (WE[5]), .\WE[6] (WE[6]), .\WE[7] (WE[7]), 
            .\WE[8] (WE[8]), .\WE[9] (WE[9]), .\WE[10] (WE[10]), .\WE[11] (WE[11]), 
            .\WE[12] (WE[12]), .\WE[13] (WE[13]), .\WE[14] (WE[14]), .\WE[15] (WE[15]), 
            .\WE[16] (WE[16]), .\WE[17] (WE[17]), .\WE[18] (WE[18]), .\WE[19] (WE[19]), 
            .\WE[20] (WE[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(359[14:22])
    \WS2812(48000000,"111111111")_U30  WS2812_18 (.sclk_c(sclk_c), .\port_status[18] (port_status[18]), 
            .ws2813_out_c_18(ws2813_out_c_18), .\Q[18] ({\Q[18] }), .\RdAddress[18] ({\RdAddress[18] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(333[13:19])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    \WS2812(48000000,"111111111")_U29  WS2812_19 (.sclk_c(sclk_c), .\port_status[19] (port_status[19]), 
            .ws2813_out_c_19(ws2813_out_c_19), .\Q[19] ({\Q[19] }), .\RdAddress[19] ({\RdAddress[19] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(344[13:19])
    \spi_slave(8,'0','0','0')  spi_port (.rx_data_cnt({Open_0, Open_1, Open_2, 
            Open_3, Open_4, rx_data_cnt[0]}), .SCLK_SLAVE_c(SCLK_SLAVE_c), 
            .rx_data_cnt_5__N_63(rx_data_cnt_5__N_63), .n50005(n50005), 
            .sclk_c(sclk_c), .RX_RDY(RX_RDY), .DATA_OUT({DATA_OUT}), .MOSI_SLAVE_c(MOSI_SLAVE_c), 
            .CSn(CSn), .CSn_SLAVE_c(CSn_SLAVE_c), .SCLK_SLAVE_c_enable_5(SCLK_SLAVE_c_enable_5));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(123[12:21])
    \WS2812(48000000,"111111111")_U33  WS2812_15 (.sclk_c(sclk_c), .\port_status[15] (port_status[15]), 
            .ws2813_out_c_15(ws2813_out_c_15), .\Q[15] ({\Q[15] }), .\RdAddress[15] ({\RdAddress[15] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(300[13:19])
    \WS2812(48000000,"111111111")_U31  WS2812_17 (.sclk_c(sclk_c), .\port_status[17] (port_status[17]), 
            .ws2813_out_c_17(ws2813_out_c_17), .\Q[17] ({\Q[17] }), .\RdAddress[17] ({\RdAddress[17] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(322[13:19])
    \WS2812(48000000,"111111111")_U26  WS2812_2 (.sclk_c(sclk_c), .\port_status[2] (port_status[2]), 
            .ws2813_out_c_2(ws2813_out_c_2), .GND_net(GND_net), .\Q[2] ({\Q[2] }), 
            .\RdAddress[2] ({\RdAddress[2] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(157[12:18])
    \WS2812(48000000,"111111111")_U36  WS2812_12 (.sclk_c(sclk_c), .\port_status[12] (port_status[12]), 
            .ws2813_out_c_12(ws2813_out_c_12), .GND_net(GND_net), .\Q[12] ({\Q[12] }), 
            .\RdAddress[12] ({\RdAddress[12] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(267[13:19])
    \WS2812(48000000,"111111111")_U23  WS2812_5 (.sclk_c(sclk_c), .\port_status[5] (port_status[5]), 
            .ws2813_out_c_5(ws2813_out_c_5), .GND_net(GND_net), .\Q[5] ({\Q[5] }), 
            .\RdAddress[5] ({\RdAddress[5] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(190[12:18])
    \WS2812(48000000,"111111111")_U24  WS2812_4 (.sclk_c(sclk_c), .\port_status[4] (port_status[4]), 
            .ws2813_out_c_4(ws2813_out_c_4), .\Q[4] ({\Q[4] }), .\RdAddress[4] ({\RdAddress[4] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(179[12:18])
    \WS2812(48000000,"111111111")_U20  WS2812_8 (.GND_net(GND_net), .sclk_c(sclk_c), 
            .\port_status[8] (port_status[8]), .ws2813_out_c_8(ws2813_out_c_8), 
            .\Q[8] ({\Q[8] }), .\RdAddress[8] ({\RdAddress[8] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(223[12:18])
    GSR GSR_INST (.GSR(n34568));
    frame_buffer_0 framebuffer9 (.WrAddress({WrAddress}), .\RdAddress[9] ({\RdAddress[9] }), 
            .Data({Data}), .\WE[9] (WE[9]), .sclk_c(sclk_c), .VCC_net(VCC_net), 
            .GND_net(GND_net), .\Q[9] ({\Q[9] })) /* synthesis NGD_DRC_MASK=1 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(229[16:30])
    \WS2812(48000000,"111111111")_U25  WS2812_3 (.sclk_c(sclk_c), .\port_status[3] (port_status[3]), 
            .ws2813_out_c_3(ws2813_out_c_3), .state({state_adj_1050}), .n13101(n13101), 
            .\Q[3] ({\Q[3] }), .\RdAddress[3] ({\RdAddress[3] }), .n41629(n41629), 
            .n10470(n10470), .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(168[12:18])
    \WS2812(48000000,"111111111")_U22  WS2812_6 (.sclk_c(sclk_c), .\port_status[6] (port_status[6]), 
            .ws2813_out_c_6(ws2813_out_c_6), .\Q[6] ({\Q[6] }), .\RdAddress[6] ({\RdAddress[6] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(201[12:18])
    \WS2812(48000000,"111111111")_U39  WS2812_0 (.\port_status[0] (port_status[0]), 
            .sclk_c(sclk_c), .ws2813_out_c_0(ws2813_out_c_0), .GND_net(GND_net), 
            .\Q[0] ({\Q[0] }), .\RdAddress[0] ({\RdAddress[0] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(135[12:18])
    \WS2812(48000000,"111111111")_U28  WS2812_1 (.sclk_c(sclk_c), .GND_net(GND_net), 
            .\port_status[1] (port_status[1]), .ws2813_out_c_1(ws2813_out_c_1), 
            .\Q[1] ({\Q[1] }), .\RdAddress[1] ({\RdAddress[1] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(146[12:18])
    \WS2812(48000000,"111111111")_U32  WS2812_16 (.sclk_c(sclk_c), .\port_status[16] (port_status[16]), 
            .ws2813_out_c_16(ws2813_out_c_16), .\Q[16] ({\Q[16] }), .\RdAddress[16] ({\RdAddress[16] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(311[13:19])
    \WS2812(48000000,"111111111")_U27  WS2812_20 (.sclk_c(sclk_c), .\port_status[20] (port_status[20]), 
            .ws2813_out_c_20(ws2813_out_c_20), .\Q[20] ({\Q[20] }), .\RdAddress[20] ({\RdAddress[20] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(355[13:19])
    \WS2812(48000000,"111111111")_U34  WS2812_14 (.GND_net(GND_net), .sclk_c(sclk_c), 
            .\port_status[14] (port_status[14]), .ws2813_out_c_14(ws2813_out_c_14), 
            .\Q[14] ({\Q[14] }), .\RdAddress[14] ({\RdAddress[14] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(289[13:19])
    \WS2812(48000000,"111111111")_U37  WS2812_11 (.GND_net(GND_net), .sclk_c(sclk_c), 
            .\port_status[11] (port_status[11]), .ws2813_out_c_11(ws2813_out_c_11), 
            .state({state_adj_1482}), .n54591(n54591), .\Q[11] ({\Q[11] }), 
            .\RdAddress[11] ({\RdAddress[11] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(256[13:19])
    \WS2812(48000000,"111111111")_U38  WS2812_10 (.sclk_c(sclk_c), .\port_status[10] (port_status[10]), 
            .ws2813_out_c_10(ws2813_out_c_10), .GND_net(GND_net), .\Q[10] ({\Q[10] }), 
            .\RdAddress[10] ({\RdAddress[10] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(245[13:19])
    \WS2812(48000000,"111111111")_U35  WS2812_13 (.sclk_c(sclk_c), .\port_status[13] (port_status[13]), 
            .ws2813_out_c_13(ws2813_out_c_13), .state({state_adj_1590}), 
            .n54583(n54583), .\Q[13] ({\Q[13] }), .\RdAddress[13] ({\RdAddress[13] }), 
            .GND_net(GND_net));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(278[13:19])
    \WS2812(48000000,"111111111")_U21  WS2812_7 (.\RdAddress[7] ({\RdAddress[7] }), 
            .sclk_c(sclk_c), .\port_status[7] (port_status[7]), .ws2813_out_c_7(ws2813_out_c_7), 
            .GND_net(GND_net), .\Q[7] ({\Q[7] }));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(212[12:18])
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111") 
//

module \WS2812(48000000,"111111111")  (sclk_c, \port_status[9] , ws2813_out_c_9, 
            GND_net, \Q[9] , \RdAddress[9] );
    input sclk_c;
    output \port_status[9] ;
    output ws2813_out_c_9;
    input GND_net;
    input [23:0]\Q[9] ;
    output [8:0]\RdAddress[9] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_2504, n35415;
    wire [31:0]n447;
    
    wire n35411, n54976, n55007;
    wire [31:0]n8212;
    
    wire sclk_c_enable_86, n54800, sclk_c_enable_87, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_90;
    wire [2:0]state_2__N_104;
    
    wire n53064, n53065;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53068, n53066, n53067, n53069, n13521, n9090, n54975, 
        n54974, n38816, n13486, n54656, n54598, n54698, n103, 
        n55006, n55005, serial_N_437, n54842;
    wire [31:0]n8036;
    
    wire n53303, n53304, n53305, n76, n48274;
    wire [31:0]bit_counter_31__N_204;
    
    wire sclk_c_enable_2323;
    wire [6:0]n15049;
    
    wire n54714;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n35593;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_2290;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_2354;
    wire [31:0]bit_counter_31__N_172;
    
    wire n48273, n48272, n48271, n53056, n53057, n53058, n53059, 
        n48270, n53060, n53061, n53062, n53063, n48269, n48268, 
        n48267, n48266, n48265, n48264, n48263;
    wire [8:0]n118;
    
    wire n48262, n38803, n48261, n1, n1_adj_925, n53302, n53301, 
        n53300, n53299, n48260, n54633, n8211, n48259, n69, n52730, 
        n15, n14, n53070, n47771, n47770, n47769, n47768, n47767, 
        n47766, n47765, n47764, n47763, n47762, n47761, n47760, 
        n47759, n47758, n47757, n47756, n47754, n47753, n47752, 
        n47751, n48449, n48448, n48447, n48446, n48445, n48444, 
        n48443, n48442, n48441, n48440, n48439, n48438, n48437, 
        n48436, n48435, n48434, n48433, n48432, n48431, n48430, 
        n48429, n48428, n48427, n48426, n48425, n48424, n48423, 
        n48422, n48421, n48420, n48419, n48418, n68, n54571, n4;
    
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2504), .CD(n35415), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2504), .CD(n35415), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54976), .SP(sclk_c_enable_2504), .CD(n35411), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n55007), .SP(sclk_c_enable_2504), .CD(n35411), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i0 (.D(n8212[0]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54800), .SP(sclk_c_enable_86), .CK(sclk_c), 
            .Q(\port_status[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_87), .CK(sclk_c), 
            .Q(ws2813_out_c_9)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_90), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_90), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_90), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    L6MUX21 i37862 (.D0(n53064), .D1(n53065), .SD(bit_counter[2]), .Z(n53068));
    L6MUX21 i37863 (.D0(n53066), .D1(n53067), .SD(bit_counter[2]), .Z(n53069));
    LUT4 i38451_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13521), .Z(sclk_c_enable_90)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38451_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13521), .Z(n9090)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 mux_2354_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13521), .Z(n54975)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2354_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2354_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13521), .Z(n54974)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2354_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 i37689_2_lut_rep_653 (.A(n38816), .B(n13486), .Z(n54656)) /* synthesis lut_function=(A (B)) */ ;
    defparam i37689_2_lut_rep_653.init = 16'h8888;
    LUT4 i1_2_lut_rep_595_3_lut (.A(n38816), .B(n13486), .C(state[1]), 
         .Z(n54598)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_595_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n38816), .B(n13486), .C(n54698), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2354_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13521), .Z(n55006)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2354_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2354_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13486), .Z(n55005)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2354_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i21986_1_lut_rep_797 (.A(state[2]), .Z(n54800)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i21986_1_lut_rep_797.init = 16'h5555;
    LUT4 i28814_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28814_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_3_lut_4_lut (.A(n54598), .B(n54842), .C(n447[7]), .D(n54698), 
         .Z(n8036[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_885 (.A(n54598), .B(n54842), .C(n447[8]), 
         .D(n54698), .Z(n8036[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_885.init = 16'hf888;
    L6MUX21 i38099 (.D0(n53303), .D1(n53304), .SD(bit_counter[2]), .Z(n53305));
    LUT4 i1_3_lut_4_lut_adj_886 (.A(n54598), .B(n54842), .C(n447[9]), 
         .D(n54698), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_886.init = 16'hf888;
    CCU2D add_3120_33 (.A0(bit_counter[31]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48274), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_33.INIT0 = 16'h5999;
    defparam add_3120_33.INIT1 = 16'h0000;
    defparam add_3120_33.INJECT1_0 = "NO";
    defparam add_3120_33.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13521), 
         .Z(sclk_c_enable_87)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_3_lut_rep_730_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_2323)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_730_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n15049[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_711_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54714)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_711_3_lut.init = 16'hf8f8;
    FD1P3AX delay_counter_i0_i1 (.D(n8212[1]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n8212[3]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n8212[7]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n8212[8]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n8212[9]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n8212[12]), .SP(sclk_c_enable_2504), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3IX pixel_i0 (.D(\Q[9] [0]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    LUT4 i38394_2_lut_rep_825 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_2354)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38394_2_lut_rep_825.init = 16'h9999;
    LUT4 i23352_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35593)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23352_2_lut_2_lut.init = 16'h8888;
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 mux_2566_i2_4_lut_4_lut (.A(n54714), .B(n54698), .C(n9090), .D(n13486), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2566_i2_4_lut_4_lut.init = 16'h5053;
    CCU2D add_3120_31 (.A0(bit_counter[29]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48273), .COUT(n48274), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_31.INIT0 = 16'h5999;
    defparam add_3120_31.INIT1 = 16'h5999;
    defparam add_3120_31.INJECT1_0 = "NO";
    defparam add_3120_31.INJECT1_1 = "NO";
    CCU2D add_3120_29 (.A0(bit_counter[27]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48272), .COUT(n48273), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_29.INIT0 = 16'h5999;
    defparam add_3120_29.INIT1 = 16'h5999;
    defparam add_3120_29.INJECT1_0 = "NO";
    defparam add_3120_29.INJECT1_1 = "NO";
    CCU2D add_3120_27 (.A0(bit_counter[25]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48271), .COUT(n48272), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_27.INIT0 = 16'h5999;
    defparam add_3120_27.INIT1 = 16'h5999;
    defparam add_3120_27.INJECT1_0 = "NO";
    defparam add_3120_27.INJECT1_1 = "NO";
    PFUMX i37858 (.BLUT(n53056), .ALUT(n53057), .C0(bit_counter[1]), .Z(n53064));
    PFUMX i37859 (.BLUT(n53058), .ALUT(n53059), .C0(bit_counter[1]), .Z(n53065));
    CCU2D add_3120_25 (.A0(bit_counter[23]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48270), .COUT(n48271), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_25.INIT0 = 16'h5999;
    defparam add_3120_25.INIT1 = 16'h5999;
    defparam add_3120_25.INJECT1_0 = "NO";
    defparam add_3120_25.INJECT1_1 = "NO";
    PFUMX i37860 (.BLUT(n53060), .ALUT(n53061), .C0(bit_counter[1]), .Z(n53066));
    PFUMX i37861 (.BLUT(n53062), .ALUT(n53063), .C0(bit_counter[1]), .Z(n53067));
    CCU2D add_3120_23 (.A0(bit_counter[21]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48269), .COUT(n48270), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_23.INIT0 = 16'h5999;
    defparam add_3120_23.INIT1 = 16'h5999;
    defparam add_3120_23.INJECT1_0 = "NO";
    defparam add_3120_23.INJECT1_1 = "NO";
    CCU2D add_3120_21 (.A0(bit_counter[19]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48268), .COUT(n48269), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_21.INIT0 = 16'h5999;
    defparam add_3120_21.INIT1 = 16'h5999;
    defparam add_3120_21.INJECT1_0 = "NO";
    defparam add_3120_21.INJECT1_1 = "NO";
    CCU2D add_3120_19 (.A0(bit_counter[17]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48267), .COUT(n48268), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_19.INIT0 = 16'h5999;
    defparam add_3120_19.INIT1 = 16'h5999;
    defparam add_3120_19.INJECT1_0 = "NO";
    defparam add_3120_19.INJECT1_1 = "NO";
    CCU2D add_3120_17 (.A0(bit_counter[15]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48266), .COUT(n48267), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_17.INIT0 = 16'h5999;
    defparam add_3120_17.INIT1 = 16'h5999;
    defparam add_3120_17.INJECT1_0 = "NO";
    defparam add_3120_17.INJECT1_1 = "NO";
    CCU2D add_3120_15 (.A0(bit_counter[13]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48265), .COUT(n48266), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_15.INIT0 = 16'h5999;
    defparam add_3120_15.INIT1 = 16'h5999;
    defparam add_3120_15.INJECT1_0 = "NO";
    defparam add_3120_15.INJECT1_1 = "NO";
    CCU2D add_3120_13 (.A0(bit_counter[11]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48264), .COUT(n48265), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_13.INIT0 = 16'h5999;
    defparam add_3120_13.INIT1 = 16'h5999;
    defparam add_3120_13.INJECT1_0 = "NO";
    defparam add_3120_13.INJECT1_1 = "NO";
    CCU2D add_3120_11 (.A0(bit_counter[9]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48263), .COUT(n48264), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_11.INIT0 = 16'h5999;
    defparam add_3120_11.INIT1 = 16'h5999;
    defparam add_3120_11.INJECT1_0 = "NO";
    defparam add_3120_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_887 (.A(state[2]), .B(n38816), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_887.init = 16'h1010;
    CCU2D add_3120_9 (.A0(bit_counter[7]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48262), .COUT(n48263), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_9.INIT0 = 16'h5999;
    defparam add_3120_9.INIT1 = 16'h5999;
    defparam add_3120_9.INJECT1_0 = "NO";
    defparam add_3120_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_888 (.A(state[2]), .B(n38816), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_888.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_889 (.A(state[2]), .B(n38816), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_889.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_890 (.A(state[2]), .B(n38816), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_890.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_891 (.A(state[2]), .B(n38816), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_891.init = 16'h1010;
    LUT4 i1_2_lut_rep_839 (.A(state[2]), .B(state[0]), .Z(n54842)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_839.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13486), 
         .D(state[1]), .Z(n38803)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13486), 
         .D(state[1]), .Z(sclk_c_enable_2290)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_3_lut_adj_892 (.A(state[2]), .B(n38816), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_892.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_893 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_893.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_894 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_894.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_895 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_895.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_896 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_896.init = 16'h4040;
    CCU2D add_3120_7 (.A0(bit_counter[5]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48261), .COUT(n48262), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_7.INIT0 = 16'h5999;
    defparam add_3120_7.INIT1 = 16'h5999;
    defparam add_3120_7.INJECT1_0 = "NO";
    defparam add_3120_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_897 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_897.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_898 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_898.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_899 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_899.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_900 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_900.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_901 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_901.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_902 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_902.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_903 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_903.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_904 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_904.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_905 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_905.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_906 (.A(state[2]), .B(n38816), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_906.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_907 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_907.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_908 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_908.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_909 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_909.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_910 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_910.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_911 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_911.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_912 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_912.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_913 (.A(state[2]), .B(n38816), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_913.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_914 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_914.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_915 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_915.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_916 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_916.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_917 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_917.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_918 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_918.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_919 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_919.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_920 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_920.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_921 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_921.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_922 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_922.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_923 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_923.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_924 (.A(state[2]), .B(n38816), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_924.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_925 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_925.init = 16'h4040;
    LUT4 i28774_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28774_2_lut.init = 16'hbbbb;
    LUT4 i28773_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_925)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28773_2_lut.init = 16'hbbbb;
    LUT4 i38096_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38096_3_lut.init = 16'hcaca;
    LUT4 i38095_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38095_3_lut.init = 16'hcaca;
    LUT4 i38094_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38094_3_lut.init = 16'hcaca;
    LUT4 i38093_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38093_3_lut.init = 16'hcaca;
    CCU2D add_3120_5 (.A0(bit_counter[3]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48260), .COUT(n48261), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_5.INIT0 = 16'h5999;
    defparam add_3120_5.INIT1 = 16'h5999;
    defparam add_3120_5.INJECT1_0 = "NO";
    defparam add_3120_5.INJECT1_1 = "NO";
    LUT4 i23199_2_lut_4_lut (.A(n54633), .B(state[0]), .C(state[1]), .D(n8211), 
         .Z(n35411)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23199_2_lut_4_lut.init = 16'hfd00;
    CCU2D add_3120_3 (.A0(bit_counter[1]), .B0(n13486), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13486), .C1(GND_net), 
          .D1(GND_net), .CIN(n48259), .COUT(n48260), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_3.INIT0 = 16'h5999;
    defparam add_3120_3.INIT1 = 16'h5999;
    defparam add_3120_3.INJECT1_0 = "NO";
    defparam add_3120_3.INJECT1_1 = "NO";
    CCU2D add_3120_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13486), .C1(GND_net), .D1(GND_net), 
          .COUT(n48259), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3120_1.INIT0 = 16'hF000;
    defparam add_3120_1.INIT1 = 16'h5999;
    defparam add_3120_1.INJECT1_0 = "NO";
    defparam add_3120_1.INJECT1_1 = "NO";
    LUT4 mux_2364_i1_4_lut (.A(n69), .B(n15049[0]), .C(n8211), .D(n52730), 
         .Z(n8212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i1_4_lut.init = 16'hcfca;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[3]), .C(n14), .D(cur_pixel[6]), 
         .Z(n38816)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    L6MUX21 i37864 (.D0(n53068), .D1(n53069), .SD(bit_counter[3]), .Z(n53070));
    LUT4 i6_4_lut (.A(cur_pixel[4]), .B(cur_pixel[2]), .C(cur_pixel[8]), 
         .D(cur_pixel[7]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47771), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47770), .COUT(n47771), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54842), .B(state[1]), .C(n54656), .D(n54633), 
         .Z(n52730)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47769), .COUT(n47770), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    LUT4 i37857_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37857_3_lut.init = 16'hcaca;
    LUT4 i37856_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37856_3_lut.init = 16'hcaca;
    LUT4 i37855_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37855_3_lut.init = 16'hcaca;
    LUT4 i37854_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37854_3_lut.init = 16'hcaca;
    LUT4 i37853_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37853_3_lut.init = 16'hcaca;
    LUT4 i37852_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37852_3_lut.init = 16'hcaca;
    LUT4 i37851_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37851_3_lut.init = 16'hcaca;
    LUT4 i37850_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37850_3_lut.init = 16'hcaca;
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47768), .COUT(n47769), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47767), .COUT(n47768), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47766), .COUT(n47767), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_86)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    PFUMX i38097 (.BLUT(n53299), .ALUT(n53300), .C0(bit_counter[1]), .Z(n53303));
    PFUMX i38098 (.BLUT(n53301), .ALUT(n53302), .C0(bit_counter[1]), .Z(n53304));
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47765), .COUT(n47766), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47764), .COUT(n47765), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47763), .COUT(n47764), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47762), .COUT(n47763), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53070), .B(n53305), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47761), .COUT(n47762), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47760), .COUT(n47761), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47759), .COUT(n47760), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 mux_2566_i1_4_lut (.A(n54656), .B(n54714), .C(n9090), .D(n54698), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2566_i1_4_lut.init = 16'h3f3a;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47758), .COUT(n47759), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47757), .COUT(n47758), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47756), .COUT(n47757), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47756), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47754), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47753), .COUT(n47754), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47752), .COUT(n47753), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    LUT4 i5_3_lut (.A(cur_pixel[5]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54656), .C(n13521), .D(n54842), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47751), .COUT(n47752), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47751), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_33916_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48449), 
          .S0(n13521));
    defparam add_33916_cout.INIT0 = 16'h0000;
    defparam add_33916_cout.INIT1 = 16'h0000;
    defparam add_33916_cout.INJECT1_0 = "NO";
    defparam add_33916_cout.INJECT1_1 = "NO";
    CCU2D add_33916_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48448), .COUT(n48449));
    defparam add_33916_31.INIT0 = 16'hf555;
    defparam add_33916_31.INIT1 = 16'h5555;
    defparam add_33916_31.INJECT1_0 = "NO";
    defparam add_33916_31.INJECT1_1 = "NO";
    CCU2D add_33916_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48447), .COUT(n48448));
    defparam add_33916_29.INIT0 = 16'hf555;
    defparam add_33916_29.INIT1 = 16'hf555;
    defparam add_33916_29.INJECT1_0 = "NO";
    defparam add_33916_29.INJECT1_1 = "NO";
    CCU2D add_33916_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48446), .COUT(n48447));
    defparam add_33916_27.INIT0 = 16'hf555;
    defparam add_33916_27.INIT1 = 16'hf555;
    defparam add_33916_27.INJECT1_0 = "NO";
    defparam add_33916_27.INJECT1_1 = "NO";
    CCU2D add_33916_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48445), .COUT(n48446));
    defparam add_33916_25.INIT0 = 16'hf555;
    defparam add_33916_25.INIT1 = 16'hf555;
    defparam add_33916_25.INJECT1_0 = "NO";
    defparam add_33916_25.INJECT1_1 = "NO";
    CCU2D add_33916_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48444), .COUT(n48445));
    defparam add_33916_23.INIT0 = 16'hf555;
    defparam add_33916_23.INIT1 = 16'hf555;
    defparam add_33916_23.INJECT1_0 = "NO";
    defparam add_33916_23.INJECT1_1 = "NO";
    CCU2D add_33916_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48443), .COUT(n48444));
    defparam add_33916_21.INIT0 = 16'hf555;
    defparam add_33916_21.INIT1 = 16'hf555;
    defparam add_33916_21.INJECT1_0 = "NO";
    defparam add_33916_21.INJECT1_1 = "NO";
    CCU2D add_33916_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48442), .COUT(n48443));
    defparam add_33916_19.INIT0 = 16'hf555;
    defparam add_33916_19.INIT1 = 16'hf555;
    defparam add_33916_19.INJECT1_0 = "NO";
    defparam add_33916_19.INJECT1_1 = "NO";
    CCU2D add_33916_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48441), .COUT(n48442));
    defparam add_33916_17.INIT0 = 16'hf555;
    defparam add_33916_17.INIT1 = 16'hf555;
    defparam add_33916_17.INJECT1_0 = "NO";
    defparam add_33916_17.INJECT1_1 = "NO";
    CCU2D add_33916_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48440), .COUT(n48441));
    defparam add_33916_15.INIT0 = 16'hf555;
    defparam add_33916_15.INIT1 = 16'hf555;
    defparam add_33916_15.INJECT1_0 = "NO";
    defparam add_33916_15.INJECT1_1 = "NO";
    CCU2D add_33916_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48439), .COUT(n48440));
    defparam add_33916_13.INIT0 = 16'hf555;
    defparam add_33916_13.INIT1 = 16'hf555;
    defparam add_33916_13.INJECT1_0 = "NO";
    defparam add_33916_13.INJECT1_1 = "NO";
    CCU2D add_33916_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48438), .COUT(n48439));
    defparam add_33916_11.INIT0 = 16'hf555;
    defparam add_33916_11.INIT1 = 16'hf555;
    defparam add_33916_11.INJECT1_0 = "NO";
    defparam add_33916_11.INJECT1_1 = "NO";
    CCU2D add_33916_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48437), .COUT(n48438));
    defparam add_33916_9.INIT0 = 16'hf555;
    defparam add_33916_9.INIT1 = 16'hf555;
    defparam add_33916_9.INJECT1_0 = "NO";
    defparam add_33916_9.INJECT1_1 = "NO";
    CCU2D add_33916_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48436), .COUT(n48437));
    defparam add_33916_7.INIT0 = 16'hf555;
    defparam add_33916_7.INIT1 = 16'hf555;
    defparam add_33916_7.INJECT1_0 = "NO";
    defparam add_33916_7.INJECT1_1 = "NO";
    CCU2D add_33916_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48435), .COUT(n48436));
    defparam add_33916_5.INIT0 = 16'hf555;
    defparam add_33916_5.INIT1 = 16'hf555;
    defparam add_33916_5.INJECT1_0 = "NO";
    defparam add_33916_5.INJECT1_1 = "NO";
    CCU2D add_33916_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48434), .COUT(n48435));
    defparam add_33916_3.INIT0 = 16'hf555;
    defparam add_33916_3.INIT1 = 16'hf555;
    defparam add_33916_3.INJECT1_0 = "NO";
    defparam add_33916_3.INJECT1_1 = "NO";
    CCU2D add_33916_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48434));
    defparam add_33916_1.INIT0 = 16'hF000;
    defparam add_33916_1.INIT1 = 16'ha666;
    defparam add_33916_1.INJECT1_0 = "NO";
    defparam add_33916_1.INJECT1_1 = "NO";
    CCU2D add_33917_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48433), 
          .S0(n13486));
    defparam add_33917_cout.INIT0 = 16'h0000;
    defparam add_33917_cout.INIT1 = 16'h0000;
    defparam add_33917_cout.INJECT1_0 = "NO";
    defparam add_33917_cout.INJECT1_1 = "NO";
    CCU2D add_33917_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48432), .COUT(n48433));
    defparam add_33917_31.INIT0 = 16'hf555;
    defparam add_33917_31.INIT1 = 16'h5555;
    defparam add_33917_31.INJECT1_0 = "NO";
    defparam add_33917_31.INJECT1_1 = "NO";
    CCU2D add_33917_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48431), .COUT(n48432));
    defparam add_33917_29.INIT0 = 16'hf555;
    defparam add_33917_29.INIT1 = 16'hf555;
    defparam add_33917_29.INJECT1_0 = "NO";
    defparam add_33917_29.INJECT1_1 = "NO";
    CCU2D add_33917_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48430), .COUT(n48431));
    defparam add_33917_27.INIT0 = 16'hf555;
    defparam add_33917_27.INIT1 = 16'hf555;
    defparam add_33917_27.INJECT1_0 = "NO";
    defparam add_33917_27.INJECT1_1 = "NO";
    CCU2D add_33917_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48429), .COUT(n48430));
    defparam add_33917_25.INIT0 = 16'hf555;
    defparam add_33917_25.INIT1 = 16'hf555;
    defparam add_33917_25.INJECT1_0 = "NO";
    defparam add_33917_25.INJECT1_1 = "NO";
    CCU2D add_33917_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48428), .COUT(n48429));
    defparam add_33917_23.INIT0 = 16'hf555;
    defparam add_33917_23.INIT1 = 16'hf555;
    defparam add_33917_23.INJECT1_0 = "NO";
    defparam add_33917_23.INJECT1_1 = "NO";
    CCU2D add_33917_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48427), .COUT(n48428));
    defparam add_33917_21.INIT0 = 16'hf555;
    defparam add_33917_21.INIT1 = 16'hf555;
    defparam add_33917_21.INJECT1_0 = "NO";
    defparam add_33917_21.INJECT1_1 = "NO";
    CCU2D add_33917_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48426), .COUT(n48427));
    defparam add_33917_19.INIT0 = 16'hf555;
    defparam add_33917_19.INIT1 = 16'hf555;
    defparam add_33917_19.INJECT1_0 = "NO";
    defparam add_33917_19.INJECT1_1 = "NO";
    CCU2D add_33917_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48425), .COUT(n48426));
    defparam add_33917_17.INIT0 = 16'hf555;
    defparam add_33917_17.INIT1 = 16'hf555;
    defparam add_33917_17.INJECT1_0 = "NO";
    defparam add_33917_17.INJECT1_1 = "NO";
    CCU2D add_33917_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48424), .COUT(n48425));
    defparam add_33917_15.INIT0 = 16'hf555;
    defparam add_33917_15.INIT1 = 16'hf555;
    defparam add_33917_15.INJECT1_0 = "NO";
    defparam add_33917_15.INJECT1_1 = "NO";
    CCU2D add_33917_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48423), .COUT(n48424));
    defparam add_33917_13.INIT0 = 16'hf555;
    defparam add_33917_13.INIT1 = 16'hf555;
    defparam add_33917_13.INJECT1_0 = "NO";
    defparam add_33917_13.INJECT1_1 = "NO";
    CCU2D add_33917_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48422), .COUT(n48423));
    defparam add_33917_11.INIT0 = 16'hf555;
    defparam add_33917_11.INIT1 = 16'hf555;
    defparam add_33917_11.INJECT1_0 = "NO";
    defparam add_33917_11.INJECT1_1 = "NO";
    CCU2D add_33917_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48421), .COUT(n48422));
    defparam add_33917_9.INIT0 = 16'hf555;
    defparam add_33917_9.INIT1 = 16'hf555;
    defparam add_33917_9.INJECT1_0 = "NO";
    defparam add_33917_9.INJECT1_1 = "NO";
    CCU2D add_33917_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48420), .COUT(n48421));
    defparam add_33917_7.INIT0 = 16'hf555;
    defparam add_33917_7.INIT1 = 16'hf555;
    defparam add_33917_7.INJECT1_0 = "NO";
    defparam add_33917_7.INJECT1_1 = "NO";
    FD1P3IX pixel_i23 (.D(\Q[9] [23]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[9] [22]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[9] [21]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[9] [20]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[9] [19]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[9] [18]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[9] [17]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[9] [16]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[9] [15]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[9] [14]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[9] [13]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[9] [12]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[9] [11]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[9] [10]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[9] [9]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[9] [8]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[9] [7]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[9] [6]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[9] [5]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[9] [4]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[9] [3]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[9] [2]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[9] [1]), .SP(sclk_c_enable_2323), .CD(n35593), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    CCU2D add_33917_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48419), .COUT(n48420));
    defparam add_33917_5.INIT0 = 16'hf555;
    defparam add_33917_5.INIT1 = 16'hf555;
    defparam add_33917_5.INJECT1_0 = "NO";
    defparam add_33917_5.INJECT1_1 = "NO";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2290), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    CCU2D add_33917_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48418), .COUT(n48419));
    defparam add_33917_3.INIT0 = 16'hf555;
    defparam add_33917_3.INIT1 = 16'hf555;
    defparam add_33917_3.INJECT1_0 = "NO";
    defparam add_33917_3.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    CCU2D add_33917_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48418));
    defparam add_33917_1.INIT0 = 16'hF000;
    defparam add_33917_1.INIT1 = 16'ha666;
    defparam add_33917_1.INJECT1_0 = "NO";
    defparam add_33917_1.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2323), 
            .CD(n35593), .CK(sclk_c), .Q(\RdAddress[9] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_695_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54698)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_695_3_lut.init = 16'hefef;
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_2354), .CD(n35593), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_926 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_926.init = 16'he0f0;
    FD1P3IX bit_counter_i3 (.D(n1_adj_925), .SP(sclk_c_enable_2354), .CD(n35593), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_927 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_927.init = 16'he0f0;
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_2354), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 i23223_4_lut (.A(sclk_c_enable_2504), .B(n54698), .C(n8211), 
         .D(n54571), .Z(n35415)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23223_4_lut.init = 16'haaa2;
    LUT4 i2376_3_lut (.A(state[2]), .B(state[1]), .C(n13521), .Z(n8211)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2376_3_lut.init = 16'ha8a8;
    LUT4 mux_2364_i2_4_lut (.A(n68), .B(n15049[0]), .C(n8211), .D(n52730), 
         .Z(n8212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2364_i4_4_lut (.A(n38803), .B(n54714), .C(n8211), .D(n4), 
         .Z(n8212[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n38816), .B(n54571), .C(n447[3]), .D(n54698), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2364_i8_4_lut (.A(n8036[7]), .B(n54714), .C(n8211), .D(n54571), 
         .Z(n8212[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i8_4_lut.init = 16'h303a;
    LUT4 mux_2364_i9_4_lut (.A(n8036[8]), .B(n54714), .C(n8211), .D(n54571), 
         .Z(n8212[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i9_4_lut.init = 16'h303a;
    LUT4 mux_2364_i10_4_lut (.A(n76), .B(n54714), .C(n8211), .D(n54571), 
         .Z(n8212[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i10_4_lut.init = 16'h303a;
    LUT4 mux_2364_i13_4_lut (.A(n54571), .B(n54714), .C(n8211), .D(n103), 
         .Z(n8212[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2364_i13_4_lut.init = 16'h3530;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    PFUMX i38977 (.BLUT(n55005), .ALUT(n55006), .C0(state[1]), .Z(n55007));
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_630 (.A(state[2]), .B(n13521), .Z(n54633)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_630.init = 16'h4444;
    LUT4 i1_2_lut_rep_568_3_lut (.A(state[2]), .B(n13521), .C(state[1]), 
         .Z(n54571)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_568_3_lut.init = 16'h4040;
    LUT4 i38596_3_lut_rep_572_4_lut (.A(state[2]), .B(n13521), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2504)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38596_3_lut_rep_572_4_lut.init = 16'hfffb;
    PFUMX i38957 (.BLUT(n54974), .ALUT(n54975), .C0(state[0]), .Z(n54976));
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2504), 
            .CD(n35415), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=234, LSE_RLINE=234 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U9
//

module frame_buffer_0_U9 (WrAddress, \RdAddress[19] , Data, \WE[19] , 
            sclk_c, VCC_net, GND_net, \Q[19] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[19] ;
    input [23:0]Data;
    input \WE[19] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[19] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[19] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[19] [0]), .ADR5(\RdAddress[19] [1]), 
            .ADR6(\RdAddress[19] [2]), .ADR7(\RdAddress[19] [3]), .ADR8(\RdAddress[19] [4]), 
            .ADR9(\RdAddress[19] [5]), .ADR10(\RdAddress[19] [6]), .ADR11(\RdAddress[19] [7]), 
            .ADR12(\RdAddress[19] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[19] [18]), .DO10(\Q[19] [19]), .DO11(\Q[19] [20]), 
            .DO12(\Q[19] [21]), .DO13(\Q[19] [22]), .DO14(\Q[19] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(339[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[19] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[19] [0]), .ADR5(\RdAddress[19] [1]), 
            .ADR6(\RdAddress[19] [2]), .ADR7(\RdAddress[19] [3]), .ADR8(\RdAddress[19] [4]), 
            .ADR9(\RdAddress[19] [5]), .ADR10(\RdAddress[19] [6]), .ADR11(\RdAddress[19] [7]), 
            .ADR12(\RdAddress[19] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[19] [9]), .DO1(\Q[19] [10]), .DO2(\Q[19] [11]), 
            .DO3(\Q[19] [12]), .DO4(\Q[19] [13]), .DO5(\Q[19] [14]), .DO6(\Q[19] [15]), 
            .DO7(\Q[19] [16]), .DO8(\Q[19] [17]), .DO9(\Q[19] [0]), .DO10(\Q[19] [1]), 
            .DO11(\Q[19] [2]), .DO12(\Q[19] [3]), .DO13(\Q[19] [4]), .DO14(\Q[19] [5]), 
            .DO15(\Q[19] [6]), .DO16(\Q[19] [7]), .DO17(\Q[19] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=339, LSE_RLINE=339 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(339[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U7
//

module frame_buffer_0_U7 (WrAddress, \RdAddress[20] , Data, \WE[20] , 
            sclk_c, VCC_net, GND_net, \Q[20] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[20] ;
    input [23:0]Data;
    input \WE[20] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[20] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[20] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[20] [0]), .ADR5(\RdAddress[20] [1]), 
            .ADR6(\RdAddress[20] [2]), .ADR7(\RdAddress[20] [3]), .ADR8(\RdAddress[20] [4]), 
            .ADR9(\RdAddress[20] [5]), .ADR10(\RdAddress[20] [6]), .ADR11(\RdAddress[20] [7]), 
            .ADR12(\RdAddress[20] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[20] [18]), .DO10(\Q[20] [19]), .DO11(\Q[20] [20]), 
            .DO12(\Q[20] [21]), .DO13(\Q[20] [22]), .DO14(\Q[20] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=350, LSE_RLINE=350 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(350[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[20] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[20] [0]), .ADR5(\RdAddress[20] [1]), 
            .ADR6(\RdAddress[20] [2]), .ADR7(\RdAddress[20] [3]), .ADR8(\RdAddress[20] [4]), 
            .ADR9(\RdAddress[20] [5]), .ADR10(\RdAddress[20] [6]), .ADR11(\RdAddress[20] [7]), 
            .ADR12(\RdAddress[20] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[20] [9]), .DO1(\Q[20] [10]), .DO2(\Q[20] [11]), 
            .DO3(\Q[20] [12]), .DO4(\Q[20] [13]), .DO5(\Q[20] [14]), .DO6(\Q[20] [15]), 
            .DO7(\Q[20] [16]), .DO8(\Q[20] [17]), .DO9(\Q[20] [0]), .DO10(\Q[20] [1]), 
            .DO11(\Q[20] [2]), .DO12(\Q[20] [3]), .DO13(\Q[20] [4]), .DO14(\Q[20] [5]), 
            .DO15(\Q[20] [6]), .DO16(\Q[20] [7]), .DO17(\Q[20] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=350, LSE_RLINE=350 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(350[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U6
//

module frame_buffer_0_U6 (WrAddress, \RdAddress[2] , Data, \WE[2] , 
            sclk_c, VCC_net, GND_net, \Q[2] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[2] ;
    input [23:0]Data;
    input \WE[2] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[2] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[2] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[2] [0]), .ADR5(\RdAddress[2] [1]), 
            .ADR6(\RdAddress[2] [2]), .ADR7(\RdAddress[2] [3]), .ADR8(\RdAddress[2] [4]), 
            .ADR9(\RdAddress[2] [5]), .ADR10(\RdAddress[2] [6]), .ADR11(\RdAddress[2] [7]), 
            .ADR12(\RdAddress[2] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[2] [18]), .DO10(\Q[2] [19]), .DO11(\Q[2] [20]), 
            .DO12(\Q[2] [21]), .DO13(\Q[2] [22]), .DO14(\Q[2] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=152, LSE_RLINE=152 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(152[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[2] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[2] [0]), .ADR5(\RdAddress[2] [1]), 
            .ADR6(\RdAddress[2] [2]), .ADR7(\RdAddress[2] [3]), .ADR8(\RdAddress[2] [4]), 
            .ADR9(\RdAddress[2] [5]), .ADR10(\RdAddress[2] [6]), .ADR11(\RdAddress[2] [7]), 
            .ADR12(\RdAddress[2] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[2] [9]), .DO1(\Q[2] [10]), .DO2(\Q[2] [11]), 
            .DO3(\Q[2] [12]), .DO4(\Q[2] [13]), .DO5(\Q[2] [14]), .DO6(\Q[2] [15]), 
            .DO7(\Q[2] [16]), .DO8(\Q[2] [17]), .DO9(\Q[2] [0]), .DO10(\Q[2] [1]), 
            .DO11(\Q[2] [2]), .DO12(\Q[2] [3]), .DO13(\Q[2] [4]), .DO14(\Q[2] [5]), 
            .DO15(\Q[2] [6]), .DO16(\Q[2] [7]), .DO17(\Q[2] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=152, LSE_RLINE=152 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(152[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U5
//

module frame_buffer_0_U5 (WrAddress, \RdAddress[3] , Data, \WE[3] , 
            sclk_c, VCC_net, GND_net, \Q[3] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[3] ;
    input [23:0]Data;
    input \WE[3] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[3] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[3] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[3] [0]), .ADR5(\RdAddress[3] [1]), 
            .ADR6(\RdAddress[3] [2]), .ADR7(\RdAddress[3] [3]), .ADR8(\RdAddress[3] [4]), 
            .ADR9(\RdAddress[3] [5]), .ADR10(\RdAddress[3] [6]), .ADR11(\RdAddress[3] [7]), 
            .ADR12(\RdAddress[3] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[3] [18]), .DO10(\Q[3] [19]), .DO11(\Q[3] [20]), 
            .DO12(\Q[3] [21]), .DO13(\Q[3] [22]), .DO14(\Q[3] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=163, LSE_RLINE=163 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(163[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[3] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[3] [0]), .ADR5(\RdAddress[3] [1]), 
            .ADR6(\RdAddress[3] [2]), .ADR7(\RdAddress[3] [3]), .ADR8(\RdAddress[3] [4]), 
            .ADR9(\RdAddress[3] [5]), .ADR10(\RdAddress[3] [6]), .ADR11(\RdAddress[3] [7]), 
            .ADR12(\RdAddress[3] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[3] [9]), .DO1(\Q[3] [10]), .DO2(\Q[3] [11]), 
            .DO3(\Q[3] [12]), .DO4(\Q[3] [13]), .DO5(\Q[3] [14]), .DO6(\Q[3] [15]), 
            .DO7(\Q[3] [16]), .DO8(\Q[3] [17]), .DO9(\Q[3] [0]), .DO10(\Q[3] [1]), 
            .DO11(\Q[3] [2]), .DO12(\Q[3] [3]), .DO13(\Q[3] [4]), .DO14(\Q[3] [5]), 
            .DO15(\Q[3] [6]), .DO16(\Q[3] [7]), .DO17(\Q[3] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=163, LSE_RLINE=163 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(163[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U4
//

module frame_buffer_0_U4 (WrAddress, \RdAddress[4] , Data, \WE[4] , 
            sclk_c, VCC_net, GND_net, \Q[4] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[4] ;
    input [23:0]Data;
    input \WE[4] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[4] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[4] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[4] [0]), .ADR5(\RdAddress[4] [1]), 
            .ADR6(\RdAddress[4] [2]), .ADR7(\RdAddress[4] [3]), .ADR8(\RdAddress[4] [4]), 
            .ADR9(\RdAddress[4] [5]), .ADR10(\RdAddress[4] [6]), .ADR11(\RdAddress[4] [7]), 
            .ADR12(\RdAddress[4] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[4] [18]), .DO10(\Q[4] [19]), .DO11(\Q[4] [20]), 
            .DO12(\Q[4] [21]), .DO13(\Q[4] [22]), .DO14(\Q[4] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=174, LSE_RLINE=174 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(174[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[4] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[4] [0]), .ADR5(\RdAddress[4] [1]), 
            .ADR6(\RdAddress[4] [2]), .ADR7(\RdAddress[4] [3]), .ADR8(\RdAddress[4] [4]), 
            .ADR9(\RdAddress[4] [5]), .ADR10(\RdAddress[4] [6]), .ADR11(\RdAddress[4] [7]), 
            .ADR12(\RdAddress[4] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[4] [9]), .DO1(\Q[4] [10]), .DO2(\Q[4] [11]), 
            .DO3(\Q[4] [12]), .DO4(\Q[4] [13]), .DO5(\Q[4] [14]), .DO6(\Q[4] [15]), 
            .DO7(\Q[4] [16]), .DO8(\Q[4] [17]), .DO9(\Q[4] [0]), .DO10(\Q[4] [1]), 
            .DO11(\Q[4] [2]), .DO12(\Q[4] [3]), .DO13(\Q[4] [4]), .DO14(\Q[4] [5]), 
            .DO15(\Q[4] [6]), .DO16(\Q[4] [7]), .DO17(\Q[4] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=174, LSE_RLINE=174 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(174[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U3
//

module frame_buffer_0_U3 (WrAddress, \RdAddress[5] , Data, \WE[5] , 
            sclk_c, VCC_net, GND_net, \Q[5] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[5] ;
    input [23:0]Data;
    input \WE[5] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[5] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[5] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[5] [0]), .ADR5(\RdAddress[5] [1]), 
            .ADR6(\RdAddress[5] [2]), .ADR7(\RdAddress[5] [3]), .ADR8(\RdAddress[5] [4]), 
            .ADR9(\RdAddress[5] [5]), .ADR10(\RdAddress[5] [6]), .ADR11(\RdAddress[5] [7]), 
            .ADR12(\RdAddress[5] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[5] [18]), .DO10(\Q[5] [19]), .DO11(\Q[5] [20]), 
            .DO12(\Q[5] [21]), .DO13(\Q[5] [22]), .DO14(\Q[5] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=185, LSE_RLINE=185 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(185[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[5] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[5] [0]), .ADR5(\RdAddress[5] [1]), 
            .ADR6(\RdAddress[5] [2]), .ADR7(\RdAddress[5] [3]), .ADR8(\RdAddress[5] [4]), 
            .ADR9(\RdAddress[5] [5]), .ADR10(\RdAddress[5] [6]), .ADR11(\RdAddress[5] [7]), 
            .ADR12(\RdAddress[5] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[5] [9]), .DO1(\Q[5] [10]), .DO2(\Q[5] [11]), 
            .DO3(\Q[5] [12]), .DO4(\Q[5] [13]), .DO5(\Q[5] [14]), .DO6(\Q[5] [15]), 
            .DO7(\Q[5] [16]), .DO8(\Q[5] [17]), .DO9(\Q[5] [0]), .DO10(\Q[5] [1]), 
            .DO11(\Q[5] [2]), .DO12(\Q[5] [3]), .DO13(\Q[5] [4]), .DO14(\Q[5] [5]), 
            .DO15(\Q[5] [6]), .DO16(\Q[5] [7]), .DO17(\Q[5] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=185, LSE_RLINE=185 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(185[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U2
//

module frame_buffer_0_U2 (WrAddress, \RdAddress[6] , Data, \WE[6] , 
            sclk_c, VCC_net, GND_net, \Q[6] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[6] ;
    input [23:0]Data;
    input \WE[6] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[6] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[6] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[6] [0]), .ADR5(\RdAddress[6] [1]), 
            .ADR6(\RdAddress[6] [2]), .ADR7(\RdAddress[6] [3]), .ADR8(\RdAddress[6] [4]), 
            .ADR9(\RdAddress[6] [5]), .ADR10(\RdAddress[6] [6]), .ADR11(\RdAddress[6] [7]), 
            .ADR12(\RdAddress[6] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[6] [18]), .DO10(\Q[6] [19]), .DO11(\Q[6] [20]), 
            .DO12(\Q[6] [21]), .DO13(\Q[6] [22]), .DO14(\Q[6] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=196, LSE_RLINE=196 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(196[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[6] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[6] [0]), .ADR5(\RdAddress[6] [1]), 
            .ADR6(\RdAddress[6] [2]), .ADR7(\RdAddress[6] [3]), .ADR8(\RdAddress[6] [4]), 
            .ADR9(\RdAddress[6] [5]), .ADR10(\RdAddress[6] [6]), .ADR11(\RdAddress[6] [7]), 
            .ADR12(\RdAddress[6] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[6] [9]), .DO1(\Q[6] [10]), .DO2(\Q[6] [11]), 
            .DO3(\Q[6] [12]), .DO4(\Q[6] [13]), .DO5(\Q[6] [14]), .DO6(\Q[6] [15]), 
            .DO7(\Q[6] [16]), .DO8(\Q[6] [17]), .DO9(\Q[6] [0]), .DO10(\Q[6] [1]), 
            .DO11(\Q[6] [2]), .DO12(\Q[6] [3]), .DO13(\Q[6] [4]), .DO14(\Q[6] [5]), 
            .DO15(\Q[6] [6]), .DO16(\Q[6] [7]), .DO17(\Q[6] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=196, LSE_RLINE=196 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(196[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U1
//

module frame_buffer_0_U1 (WrAddress, \RdAddress[7] , Data, \WE[7] , 
            sclk_c, VCC_net, GND_net, \Q[7] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[7] ;
    input [23:0]Data;
    input \WE[7] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[7] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[7] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[7] [0]), .ADR5(\RdAddress[7] [1]), 
            .ADR6(\RdAddress[7] [2]), .ADR7(\RdAddress[7] [3]), .ADR8(\RdAddress[7] [4]), 
            .ADR9(\RdAddress[7] [5]), .ADR10(\RdAddress[7] [6]), .ADR11(\RdAddress[7] [7]), 
            .ADR12(\RdAddress[7] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[7] [18]), .DO10(\Q[7] [19]), .DO11(\Q[7] [20]), 
            .DO12(\Q[7] [21]), .DO13(\Q[7] [22]), .DO14(\Q[7] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=207, LSE_RLINE=207 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(207[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[7] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[7] [0]), .ADR5(\RdAddress[7] [1]), 
            .ADR6(\RdAddress[7] [2]), .ADR7(\RdAddress[7] [3]), .ADR8(\RdAddress[7] [4]), 
            .ADR9(\RdAddress[7] [5]), .ADR10(\RdAddress[7] [6]), .ADR11(\RdAddress[7] [7]), 
            .ADR12(\RdAddress[7] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[7] [9]), .DO1(\Q[7] [10]), .DO2(\Q[7] [11]), 
            .DO3(\Q[7] [12]), .DO4(\Q[7] [13]), .DO5(\Q[7] [14]), .DO6(\Q[7] [15]), 
            .DO7(\Q[7] [16]), .DO8(\Q[7] [17]), .DO9(\Q[7] [0]), .DO10(\Q[7] [1]), 
            .DO11(\Q[7] [2]), .DO12(\Q[7] [3]), .DO13(\Q[7] [4]), .DO14(\Q[7] [5]), 
            .DO15(\Q[7] [6]), .DO16(\Q[7] [7]), .DO17(\Q[7] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=207, LSE_RLINE=207 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(207[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U0
//

module frame_buffer_0_U0 (WrAddress, \RdAddress[8] , Data, \WE[8] , 
            sclk_c, VCC_net, GND_net, \Q[8] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[8] ;
    input [23:0]Data;
    input \WE[8] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[8] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[8] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[8] [0]), .ADR5(\RdAddress[8] [1]), 
            .ADR6(\RdAddress[8] [2]), .ADR7(\RdAddress[8] [3]), .ADR8(\RdAddress[8] [4]), 
            .ADR9(\RdAddress[8] [5]), .ADR10(\RdAddress[8] [6]), .ADR11(\RdAddress[8] [7]), 
            .ADR12(\RdAddress[8] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[8] [18]), .DO10(\Q[8] [19]), .DO11(\Q[8] [20]), 
            .DO12(\Q[8] [21]), .DO13(\Q[8] [22]), .DO14(\Q[8] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=218, LSE_RLINE=218 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(218[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[8] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[8] [0]), .ADR5(\RdAddress[8] [1]), 
            .ADR6(\RdAddress[8] [2]), .ADR7(\RdAddress[8] [3]), .ADR8(\RdAddress[8] [4]), 
            .ADR9(\RdAddress[8] [5]), .ADR10(\RdAddress[8] [6]), .ADR11(\RdAddress[8] [7]), 
            .ADR12(\RdAddress[8] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[8] [9]), .DO1(\Q[8] [10]), .DO2(\Q[8] [11]), 
            .DO3(\Q[8] [12]), .DO4(\Q[8] [13]), .DO5(\Q[8] [14]), .DO6(\Q[8] [15]), 
            .DO7(\Q[8] [16]), .DO8(\Q[8] [17]), .DO9(\Q[8] [0]), .DO10(\Q[8] [1]), 
            .DO11(\Q[8] [2]), .DO12(\Q[8] [3]), .DO13(\Q[8] [4]), .DO14(\Q[8] [5]), 
            .DO15(\Q[8] [6]), .DO16(\Q[8] [7]), .DO17(\Q[8] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=218, LSE_RLINE=218 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(218[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U19
//

module frame_buffer_0_U19 (WrAddress, \RdAddress[0] , Data, \WE[0] , 
            sclk_c, VCC_net, GND_net, \Q[0] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[0] ;
    input [23:0]Data;
    input \WE[0] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[0] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[0] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[0] [0]), .ADR5(\RdAddress[0] [1]), 
            .ADR6(\RdAddress[0] [2]), .ADR7(\RdAddress[0] [3]), .ADR8(\RdAddress[0] [4]), 
            .ADR9(\RdAddress[0] [5]), .ADR10(\RdAddress[0] [6]), .ADR11(\RdAddress[0] [7]), 
            .ADR12(\RdAddress[0] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[0] [18]), .DO10(\Q[0] [19]), .DO11(\Q[0] [20]), 
            .DO12(\Q[0] [21]), .DO13(\Q[0] [22]), .DO14(\Q[0] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=130, LSE_RLINE=130 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(130[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[0] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[0] [0]), .ADR5(\RdAddress[0] [1]), 
            .ADR6(\RdAddress[0] [2]), .ADR7(\RdAddress[0] [3]), .ADR8(\RdAddress[0] [4]), 
            .ADR9(\RdAddress[0] [5]), .ADR10(\RdAddress[0] [6]), .ADR11(\RdAddress[0] [7]), 
            .ADR12(\RdAddress[0] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[0] [9]), .DO1(\Q[0] [10]), .DO2(\Q[0] [11]), 
            .DO3(\Q[0] [12]), .DO4(\Q[0] [13]), .DO5(\Q[0] [14]), .DO6(\Q[0] [15]), 
            .DO7(\Q[0] [16]), .DO8(\Q[0] [17]), .DO9(\Q[0] [0]), .DO10(\Q[0] [1]), 
            .DO11(\Q[0] [2]), .DO12(\Q[0] [3]), .DO13(\Q[0] [4]), .DO14(\Q[0] [5]), 
            .DO15(\Q[0] [6]), .DO16(\Q[0] [7]), .DO17(\Q[0] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=130, LSE_RLINE=130 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(130[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U18
//

module frame_buffer_0_U18 (WrAddress, \RdAddress[10] , Data, \WE[10] , 
            sclk_c, VCC_net, GND_net, \Q[10] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[10] ;
    input [23:0]Data;
    input \WE[10] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[10] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[10] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[10] [0]), .ADR5(\RdAddress[10] [1]), 
            .ADR6(\RdAddress[10] [2]), .ADR7(\RdAddress[10] [3]), .ADR8(\RdAddress[10] [4]), 
            .ADR9(\RdAddress[10] [5]), .ADR10(\RdAddress[10] [6]), .ADR11(\RdAddress[10] [7]), 
            .ADR12(\RdAddress[10] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[10] [18]), .DO10(\Q[10] [19]), .DO11(\Q[10] [20]), 
            .DO12(\Q[10] [21]), .DO13(\Q[10] [22]), .DO14(\Q[10] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=240, LSE_RLINE=240 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(240[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[10] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[10] [0]), .ADR5(\RdAddress[10] [1]), 
            .ADR6(\RdAddress[10] [2]), .ADR7(\RdAddress[10] [3]), .ADR8(\RdAddress[10] [4]), 
            .ADR9(\RdAddress[10] [5]), .ADR10(\RdAddress[10] [6]), .ADR11(\RdAddress[10] [7]), 
            .ADR12(\RdAddress[10] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[10] [9]), .DO1(\Q[10] [10]), .DO2(\Q[10] [11]), 
            .DO3(\Q[10] [12]), .DO4(\Q[10] [13]), .DO5(\Q[10] [14]), .DO6(\Q[10] [15]), 
            .DO7(\Q[10] [16]), .DO8(\Q[10] [17]), .DO9(\Q[10] [0]), .DO10(\Q[10] [1]), 
            .DO11(\Q[10] [2]), .DO12(\Q[10] [3]), .DO13(\Q[10] [4]), .DO14(\Q[10] [5]), 
            .DO15(\Q[10] [6]), .DO16(\Q[10] [7]), .DO17(\Q[10] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=240, LSE_RLINE=240 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(240[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U17
//

module frame_buffer_0_U17 (WrAddress, \RdAddress[11] , Data, \WE[11] , 
            sclk_c, VCC_net, GND_net, \Q[11] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[11] ;
    input [23:0]Data;
    input \WE[11] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[11] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[11] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[11] [0]), .ADR5(\RdAddress[11] [1]), 
            .ADR6(\RdAddress[11] [2]), .ADR7(\RdAddress[11] [3]), .ADR8(\RdAddress[11] [4]), 
            .ADR9(\RdAddress[11] [5]), .ADR10(\RdAddress[11] [6]), .ADR11(\RdAddress[11] [7]), 
            .ADR12(\RdAddress[11] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[11] [18]), .DO10(\Q[11] [19]), .DO11(\Q[11] [20]), 
            .DO12(\Q[11] [21]), .DO13(\Q[11] [22]), .DO14(\Q[11] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=251, LSE_RLINE=251 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(251[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[11] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[11] [0]), .ADR5(\RdAddress[11] [1]), 
            .ADR6(\RdAddress[11] [2]), .ADR7(\RdAddress[11] [3]), .ADR8(\RdAddress[11] [4]), 
            .ADR9(\RdAddress[11] [5]), .ADR10(\RdAddress[11] [6]), .ADR11(\RdAddress[11] [7]), 
            .ADR12(\RdAddress[11] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[11] [9]), .DO1(\Q[11] [10]), .DO2(\Q[11] [11]), 
            .DO3(\Q[11] [12]), .DO4(\Q[11] [13]), .DO5(\Q[11] [14]), .DO6(\Q[11] [15]), 
            .DO7(\Q[11] [16]), .DO8(\Q[11] [17]), .DO9(\Q[11] [0]), .DO10(\Q[11] [1]), 
            .DO11(\Q[11] [2]), .DO12(\Q[11] [3]), .DO13(\Q[11] [4]), .DO14(\Q[11] [5]), 
            .DO15(\Q[11] [6]), .DO16(\Q[11] [7]), .DO17(\Q[11] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=251, LSE_RLINE=251 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(251[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U16
//

module frame_buffer_0_U16 (WrAddress, \RdAddress[12] , Data, \WE[12] , 
            sclk_c, VCC_net, GND_net, \Q[12] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[12] ;
    input [23:0]Data;
    input \WE[12] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[12] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[12] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[12] [0]), .ADR5(\RdAddress[12] [1]), 
            .ADR6(\RdAddress[12] [2]), .ADR7(\RdAddress[12] [3]), .ADR8(\RdAddress[12] [4]), 
            .ADR9(\RdAddress[12] [5]), .ADR10(\RdAddress[12] [6]), .ADR11(\RdAddress[12] [7]), 
            .ADR12(\RdAddress[12] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[12] [18]), .DO10(\Q[12] [19]), .DO11(\Q[12] [20]), 
            .DO12(\Q[12] [21]), .DO13(\Q[12] [22]), .DO14(\Q[12] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=262, LSE_RLINE=262 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(262[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[12] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[12] [0]), .ADR5(\RdAddress[12] [1]), 
            .ADR6(\RdAddress[12] [2]), .ADR7(\RdAddress[12] [3]), .ADR8(\RdAddress[12] [4]), 
            .ADR9(\RdAddress[12] [5]), .ADR10(\RdAddress[12] [6]), .ADR11(\RdAddress[12] [7]), 
            .ADR12(\RdAddress[12] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[12] [9]), .DO1(\Q[12] [10]), .DO2(\Q[12] [11]), 
            .DO3(\Q[12] [12]), .DO4(\Q[12] [13]), .DO5(\Q[12] [14]), .DO6(\Q[12] [15]), 
            .DO7(\Q[12] [16]), .DO8(\Q[12] [17]), .DO9(\Q[12] [0]), .DO10(\Q[12] [1]), 
            .DO11(\Q[12] [2]), .DO12(\Q[12] [3]), .DO13(\Q[12] [4]), .DO14(\Q[12] [5]), 
            .DO15(\Q[12] [6]), .DO16(\Q[12] [7]), .DO17(\Q[12] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=262, LSE_RLINE=262 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(262[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U15
//

module frame_buffer_0_U15 (WrAddress, \RdAddress[13] , Data, \WE[13] , 
            sclk_c, VCC_net, GND_net, \Q[13] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[13] ;
    input [23:0]Data;
    input \WE[13] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[13] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[13] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[13] [0]), .ADR5(\RdAddress[13] [1]), 
            .ADR6(\RdAddress[13] [2]), .ADR7(\RdAddress[13] [3]), .ADR8(\RdAddress[13] [4]), 
            .ADR9(\RdAddress[13] [5]), .ADR10(\RdAddress[13] [6]), .ADR11(\RdAddress[13] [7]), 
            .ADR12(\RdAddress[13] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[13] [18]), .DO10(\Q[13] [19]), .DO11(\Q[13] [20]), 
            .DO12(\Q[13] [21]), .DO13(\Q[13] [22]), .DO14(\Q[13] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=273, LSE_RLINE=273 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(273[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[13] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[13] [0]), .ADR5(\RdAddress[13] [1]), 
            .ADR6(\RdAddress[13] [2]), .ADR7(\RdAddress[13] [3]), .ADR8(\RdAddress[13] [4]), 
            .ADR9(\RdAddress[13] [5]), .ADR10(\RdAddress[13] [6]), .ADR11(\RdAddress[13] [7]), 
            .ADR12(\RdAddress[13] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[13] [9]), .DO1(\Q[13] [10]), .DO2(\Q[13] [11]), 
            .DO3(\Q[13] [12]), .DO4(\Q[13] [13]), .DO5(\Q[13] [14]), .DO6(\Q[13] [15]), 
            .DO7(\Q[13] [16]), .DO8(\Q[13] [17]), .DO9(\Q[13] [0]), .DO10(\Q[13] [1]), 
            .DO11(\Q[13] [2]), .DO12(\Q[13] [3]), .DO13(\Q[13] [4]), .DO14(\Q[13] [5]), 
            .DO15(\Q[13] [6]), .DO16(\Q[13] [7]), .DO17(\Q[13] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=273, LSE_RLINE=273 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(273[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U14
//

module frame_buffer_0_U14 (WrAddress, \RdAddress[14] , Data, \WE[14] , 
            sclk_c, VCC_net, GND_net, \Q[14] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[14] ;
    input [23:0]Data;
    input \WE[14] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[14] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[14] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[14] [0]), .ADR5(\RdAddress[14] [1]), 
            .ADR6(\RdAddress[14] [2]), .ADR7(\RdAddress[14] [3]), .ADR8(\RdAddress[14] [4]), 
            .ADR9(\RdAddress[14] [5]), .ADR10(\RdAddress[14] [6]), .ADR11(\RdAddress[14] [7]), 
            .ADR12(\RdAddress[14] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[14] [18]), .DO10(\Q[14] [19]), .DO11(\Q[14] [20]), 
            .DO12(\Q[14] [21]), .DO13(\Q[14] [22]), .DO14(\Q[14] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=284, LSE_RLINE=284 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(284[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[14] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[14] [0]), .ADR5(\RdAddress[14] [1]), 
            .ADR6(\RdAddress[14] [2]), .ADR7(\RdAddress[14] [3]), .ADR8(\RdAddress[14] [4]), 
            .ADR9(\RdAddress[14] [5]), .ADR10(\RdAddress[14] [6]), .ADR11(\RdAddress[14] [7]), 
            .ADR12(\RdAddress[14] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[14] [9]), .DO1(\Q[14] [10]), .DO2(\Q[14] [11]), 
            .DO3(\Q[14] [12]), .DO4(\Q[14] [13]), .DO5(\Q[14] [14]), .DO6(\Q[14] [15]), 
            .DO7(\Q[14] [16]), .DO8(\Q[14] [17]), .DO9(\Q[14] [0]), .DO10(\Q[14] [1]), 
            .DO11(\Q[14] [2]), .DO12(\Q[14] [3]), .DO13(\Q[14] [4]), .DO14(\Q[14] [5]), 
            .DO15(\Q[14] [6]), .DO16(\Q[14] [7]), .DO17(\Q[14] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=284, LSE_RLINE=284 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(284[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U13
//

module frame_buffer_0_U13 (WrAddress, \RdAddress[15] , Data, \WE[15] , 
            sclk_c, VCC_net, GND_net, \Q[15] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[15] ;
    input [23:0]Data;
    input \WE[15] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[15] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[15] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[15] [0]), .ADR5(\RdAddress[15] [1]), 
            .ADR6(\RdAddress[15] [2]), .ADR7(\RdAddress[15] [3]), .ADR8(\RdAddress[15] [4]), 
            .ADR9(\RdAddress[15] [5]), .ADR10(\RdAddress[15] [6]), .ADR11(\RdAddress[15] [7]), 
            .ADR12(\RdAddress[15] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[15] [18]), .DO10(\Q[15] [19]), .DO11(\Q[15] [20]), 
            .DO12(\Q[15] [21]), .DO13(\Q[15] [22]), .DO14(\Q[15] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=295, LSE_RLINE=295 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(295[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[15] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[15] [0]), .ADR5(\RdAddress[15] [1]), 
            .ADR6(\RdAddress[15] [2]), .ADR7(\RdAddress[15] [3]), .ADR8(\RdAddress[15] [4]), 
            .ADR9(\RdAddress[15] [5]), .ADR10(\RdAddress[15] [6]), .ADR11(\RdAddress[15] [7]), 
            .ADR12(\RdAddress[15] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[15] [9]), .DO1(\Q[15] [10]), .DO2(\Q[15] [11]), 
            .DO3(\Q[15] [12]), .DO4(\Q[15] [13]), .DO5(\Q[15] [14]), .DO6(\Q[15] [15]), 
            .DO7(\Q[15] [16]), .DO8(\Q[15] [17]), .DO9(\Q[15] [0]), .DO10(\Q[15] [1]), 
            .DO11(\Q[15] [2]), .DO12(\Q[15] [3]), .DO13(\Q[15] [4]), .DO14(\Q[15] [5]), 
            .DO15(\Q[15] [6]), .DO16(\Q[15] [7]), .DO17(\Q[15] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=295, LSE_RLINE=295 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(295[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U12
//

module frame_buffer_0_U12 (WrAddress, \RdAddress[16] , Data, \WE[16] , 
            sclk_c, VCC_net, GND_net, \Q[16] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[16] ;
    input [23:0]Data;
    input \WE[16] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[16] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[16] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[16] [0]), .ADR5(\RdAddress[16] [1]), 
            .ADR6(\RdAddress[16] [2]), .ADR7(\RdAddress[16] [3]), .ADR8(\RdAddress[16] [4]), 
            .ADR9(\RdAddress[16] [5]), .ADR10(\RdAddress[16] [6]), .ADR11(\RdAddress[16] [7]), 
            .ADR12(\RdAddress[16] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[16] [18]), .DO10(\Q[16] [19]), .DO11(\Q[16] [20]), 
            .DO12(\Q[16] [21]), .DO13(\Q[16] [22]), .DO14(\Q[16] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=306, LSE_RLINE=306 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(306[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[16] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[16] [0]), .ADR5(\RdAddress[16] [1]), 
            .ADR6(\RdAddress[16] [2]), .ADR7(\RdAddress[16] [3]), .ADR8(\RdAddress[16] [4]), 
            .ADR9(\RdAddress[16] [5]), .ADR10(\RdAddress[16] [6]), .ADR11(\RdAddress[16] [7]), 
            .ADR12(\RdAddress[16] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[16] [9]), .DO1(\Q[16] [10]), .DO2(\Q[16] [11]), 
            .DO3(\Q[16] [12]), .DO4(\Q[16] [13]), .DO5(\Q[16] [14]), .DO6(\Q[16] [15]), 
            .DO7(\Q[16] [16]), .DO8(\Q[16] [17]), .DO9(\Q[16] [0]), .DO10(\Q[16] [1]), 
            .DO11(\Q[16] [2]), .DO12(\Q[16] [3]), .DO13(\Q[16] [4]), .DO14(\Q[16] [5]), 
            .DO15(\Q[16] [6]), .DO16(\Q[16] [7]), .DO17(\Q[16] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=306, LSE_RLINE=306 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(306[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U11
//

module frame_buffer_0_U11 (WrAddress, \RdAddress[17] , Data, \WE[17] , 
            sclk_c, VCC_net, GND_net, \Q[17] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[17] ;
    input [23:0]Data;
    input \WE[17] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[17] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[17] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[17] [0]), .ADR5(\RdAddress[17] [1]), 
            .ADR6(\RdAddress[17] [2]), .ADR7(\RdAddress[17] [3]), .ADR8(\RdAddress[17] [4]), 
            .ADR9(\RdAddress[17] [5]), .ADR10(\RdAddress[17] [6]), .ADR11(\RdAddress[17] [7]), 
            .ADR12(\RdAddress[17] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[17] [18]), .DO10(\Q[17] [19]), .DO11(\Q[17] [20]), 
            .DO12(\Q[17] [21]), .DO13(\Q[17] [22]), .DO14(\Q[17] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(317[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[17] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[17] [0]), .ADR5(\RdAddress[17] [1]), 
            .ADR6(\RdAddress[17] [2]), .ADR7(\RdAddress[17] [3]), .ADR8(\RdAddress[17] [4]), 
            .ADR9(\RdAddress[17] [5]), .ADR10(\RdAddress[17] [6]), .ADR11(\RdAddress[17] [7]), 
            .ADR12(\RdAddress[17] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[17] [9]), .DO1(\Q[17] [10]), .DO2(\Q[17] [11]), 
            .DO3(\Q[17] [12]), .DO4(\Q[17] [13]), .DO5(\Q[17] [14]), .DO6(\Q[17] [15]), 
            .DO7(\Q[17] [16]), .DO8(\Q[17] [17]), .DO9(\Q[17] [0]), .DO10(\Q[17] [1]), 
            .DO11(\Q[17] [2]), .DO12(\Q[17] [3]), .DO13(\Q[17] [4]), .DO14(\Q[17] [5]), 
            .DO15(\Q[17] [6]), .DO16(\Q[17] [7]), .DO17(\Q[17] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=317, LSE_RLINE=317 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(317[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U10
//

module frame_buffer_0_U10 (WrAddress, \RdAddress[18] , Data, \WE[18] , 
            sclk_c, VCC_net, GND_net, \Q[18] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[18] ;
    input [23:0]Data;
    input \WE[18] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[18] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[18] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[18] [0]), .ADR5(\RdAddress[18] [1]), 
            .ADR6(\RdAddress[18] [2]), .ADR7(\RdAddress[18] [3]), .ADR8(\RdAddress[18] [4]), 
            .ADR9(\RdAddress[18] [5]), .ADR10(\RdAddress[18] [6]), .ADR11(\RdAddress[18] [7]), 
            .ADR12(\RdAddress[18] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[18] [18]), .DO10(\Q[18] [19]), .DO11(\Q[18] [20]), 
            .DO12(\Q[18] [21]), .DO13(\Q[18] [22]), .DO14(\Q[18] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=328, LSE_RLINE=328 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(328[17:31])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[18] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[18] [0]), .ADR5(\RdAddress[18] [1]), 
            .ADR6(\RdAddress[18] [2]), .ADR7(\RdAddress[18] [3]), .ADR8(\RdAddress[18] [4]), 
            .ADR9(\RdAddress[18] [5]), .ADR10(\RdAddress[18] [6]), .ADR11(\RdAddress[18] [7]), 
            .ADR12(\RdAddress[18] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[18] [9]), .DO1(\Q[18] [10]), .DO2(\Q[18] [11]), 
            .DO3(\Q[18] [12]), .DO4(\Q[18] [13]), .DO5(\Q[18] [14]), .DO6(\Q[18] [15]), 
            .DO7(\Q[18] [16]), .DO8(\Q[18] [17]), .DO9(\Q[18] [0]), .DO10(\Q[18] [1]), 
            .DO11(\Q[18] [2]), .DO12(\Q[18] [3]), .DO13(\Q[18] [4]), .DO14(\Q[18] [5]), 
            .DO15(\Q[18] [6]), .DO16(\Q[18] [7]), .DO17(\Q[18] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=17, LSE_RCOL=31, LSE_LLINE=328, LSE_RLINE=328 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(328[17:31])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module frame_buffer_0_U8
//

module frame_buffer_0_U8 (WrAddress, \RdAddress[1] , Data, \WE[1] , 
            sclk_c, VCC_net, GND_net, \Q[1] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[1] ;
    input [23:0]Data;
    input \WE[1] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[1] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[1] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[1] [0]), .ADR5(\RdAddress[1] [1]), 
            .ADR6(\RdAddress[1] [2]), .ADR7(\RdAddress[1] [3]), .ADR8(\RdAddress[1] [4]), 
            .ADR9(\RdAddress[1] [5]), .ADR10(\RdAddress[1] [6]), .ADR11(\RdAddress[1] [7]), 
            .ADR12(\RdAddress[1] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[1] [18]), .DO10(\Q[1] [19]), .DO11(\Q[1] [20]), 
            .DO12(\Q[1] [21]), .DO13(\Q[1] [22]), .DO14(\Q[1] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=141, LSE_RLINE=141 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(141[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[1] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[1] [0]), .ADR5(\RdAddress[1] [1]), 
            .ADR6(\RdAddress[1] [2]), .ADR7(\RdAddress[1] [3]), .ADR8(\RdAddress[1] [4]), 
            .ADR9(\RdAddress[1] [5]), .ADR10(\RdAddress[1] [6]), .ADR11(\RdAddress[1] [7]), 
            .ADR12(\RdAddress[1] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[1] [9]), .DO1(\Q[1] [10]), .DO2(\Q[1] [11]), 
            .DO3(\Q[1] [12]), .DO4(\Q[1] [13]), .DO5(\Q[1] [14]), .DO6(\Q[1] [15]), 
            .DO7(\Q[1] [16]), .DO8(\Q[1] [17]), .DO9(\Q[1] [0]), .DO10(\Q[1] [1]), 
            .DO11(\Q[1] [2]), .DO12(\Q[1] [3]), .DO13(\Q[1] [4]), .DO14(\Q[1] [5]), 
            .DO15(\Q[1] [6]), .DO16(\Q[1] [7]), .DO17(\Q[1] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=141, LSE_RLINE=141 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(141[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module \load_mem(48000000) 
//

module \load_mem(48000000)  (GND_net, Data, sclk_c, CSn, WrAddress, 
            \WE[0] , DATA_OUT, RX_RDY, \WE[1] , \WE[2] , \WE[3] , 
            \WE[4] , \WE[5] , \WE[6] , \WE[7] , \WE[8] , \WE[9] , 
            \WE[10] , \WE[11] , \WE[12] , \WE[13] , \WE[14] , \WE[15] , 
            \WE[16] , \WE[17] , \WE[18] , \WE[19] , \WE[20] );
    input GND_net;
    output [23:0]Data;
    input sclk_c;
    output CSn;
    output [8:0]WrAddress;
    output \WE[0] ;
    input [7:0]DATA_OUT;
    input RX_RDY;
    output \WE[1] ;
    output \WE[2] ;
    output \WE[3] ;
    output \WE[4] ;
    output \WE[5] ;
    output \WE[6] ;
    output \WE[7] ;
    output \WE[8] ;
    output \WE[9] ;
    output \WE[10] ;
    output \WE[11] ;
    output \WE[12] ;
    output \WE[13] ;
    output \WE[14] ;
    output \WE[15] ;
    output \WE[16] ;
    output \WE[17] ;
    output \WE[18] ;
    output \WE[19] ;
    output \WE[20] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n47550, n54553, n14326;
    wire [31:0]spi_byte_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(33[12:28])
    wire [31:0]n1337;
    
    wire n14536, n47549;
    wire [31:0]spi_byte_counter_31__N_760;
    
    wire n47548, n47547, n47546, n47545, n47544, n47543, n47542, 
        n47541, n47540, n47539, n47538, n47537, n47536, n47535, 
        sclk_c_enable_1260, sclk_c_enable_1028;
    wire [23:0]WrData_23__N_691;
    
    wire sclk_c_enable_189, SPI_CS_N_880, sclk_c_enable_1283;
    wire [8:0]WrAddr_8__N_747;
    
    wire sclk_c_enable_1315;
    wire [1:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    wire [23:0]WrEnable_23__N_824;
    wire [31:0]spi_byte_timeout;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(34[12:28])
    
    wire sclk_c_enable_224;
    wire [31:0]n1568;
    
    wire sclk_c_enable_205;
    wire [31:0]spi_byte_timeout_31__N_595;
    
    wire n55547, n48577, n14466, n48576, n48575, n48574;
    wire [31:0]index;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(35[12:17])
    
    wire n48573, n48572, n48571, n48570, n48569, n48568, n48567, 
        n48566, n48565, n15, n48564, n15_adj_916, n15_adj_917, n14501;
    wire [31:0]n869;
    
    wire n30, n48563, n55545, n98, n44072, n55544, n14571;
    wire [31:0]fb;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(30[12:14])
    
    wire n8, n8_adj_918, n8_adj_919, n8_adj_920, n8_adj_921, n48562, 
        n54678, n51598, n14361, n55003, n55002;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(32[12:25])
    
    wire sclk_c_enable_1027;
    wire [31:0]delay_counter_31__N_531;
    
    wire n54680, n36657, n1, sclk_c_enable_1092;
    wire [31:0]index_31__N_848;
    
    wire n54679, n14396, n54622, n14431, n131, n1_adj_922, n54628;
    wire [31:0]n830;
    
    wire sclk_c_enable_2505, n1_adj_923, sclk_c_enable_1111, n36653;
    wire [31:0]fb_31__N_715;
    
    wire n54742, n51592, sclk_c_enable_1268, sclk_c_enable_1276, sclk_c_enable_1284, 
        n52919, n6, n54881, n54880;
    wire [23:0]n2;
    
    wire n54741, n49273, n54681;
    wire [31:0]delay_counter_31__N_659;
    
    wire n50606, n50674, n48210, n48209, n48208, n48207, n48206, 
        n48205, n48204, n48203, n48202, n48201, n48200, n48199, 
        n48198, n48197, n48196, n49038, n49037, n49036, n49035, 
        n49034, n49033, n49032, n49031, n48195, n49030, n49029, 
        n49028, n49027, n49026, n49025, n49024, n48194, n48193, 
        n48192, n48191, n48190, n48189, n48188, n48187, n48186, 
        n48185, n48184, n48183, n48182, n48181, n48991, n48990, 
        n48989, n48988, n48987, n48986, n48985, n48984, n48983, 
        n48982, n48981, n48980, n48979, n48180, n48978, n48977, 
        n48976, n48975, n48974, n48973, n48972, n48971, n48970, 
        n48969, n48968, n48967, n48179, n48178, n48177, n48176, 
        n48175, n48174, n48173, n48966, n48172, n48171, n48170, 
        n48169, n48168, n48965, n48964, n48963, n48167, n48166, 
        n48165, n48164, n48962, n48163, n47914, n47913, n47912, 
        n47911, n47910, n47909, n47908, n47907, n47906, n47905, 
        n47904, n47903, n47902, n47901, n47900, n47899, n48417, 
        n48416, n48415, n48414, n48413, n48412, n48411, n48410, 
        n48409, n48408, n48407, n48406, n48405, n48404, n48403, 
        n48833, n48832, n48831, n48830, n48829, n48828, n48827, 
        n48826, n48825, n48824, n48823, n48822, n48821, n48820, 
        n48819, n48818, n7, n47834, n47833, n47832, n47831, n47830, 
        n47829, n47828, n47827, n47826, n47825, n47824, n47823, 
        n47822, n47821, n47820, n47819;
    
    CCU2D sub_3241_add_2_33 (.A0(n54553), .B0(n14326), .C0(spi_byte_counter[31]), 
          .D0(n1337[31]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47550), .S1(n14536));
    defparam sub_3241_add_2_33.INIT0 = 16'h078f;
    defparam sub_3241_add_2_33.INIT1 = 16'h0000;
    defparam sub_3241_add_2_33.INJECT1_0 = "NO";
    defparam sub_3241_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_31 (.A0(spi_byte_counter_31__N_760[29]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[30]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47549), .COUT(n47550));
    defparam sub_3241_add_2_31.INIT0 = 16'hf555;
    defparam sub_3241_add_2_31.INIT1 = 16'hf555;
    defparam sub_3241_add_2_31.INJECT1_0 = "NO";
    defparam sub_3241_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_29 (.A0(spi_byte_counter_31__N_760[27]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[28]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47548), .COUT(n47549));
    defparam sub_3241_add_2_29.INIT0 = 16'hf555;
    defparam sub_3241_add_2_29.INIT1 = 16'hf555;
    defparam sub_3241_add_2_29.INJECT1_0 = "NO";
    defparam sub_3241_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_27 (.A0(spi_byte_counter_31__N_760[25]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[26]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47547), .COUT(n47548));
    defparam sub_3241_add_2_27.INIT0 = 16'hf555;
    defparam sub_3241_add_2_27.INIT1 = 16'hf555;
    defparam sub_3241_add_2_27.INJECT1_0 = "NO";
    defparam sub_3241_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_25 (.A0(spi_byte_counter_31__N_760[23]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[24]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47546), .COUT(n47547));
    defparam sub_3241_add_2_25.INIT0 = 16'hf555;
    defparam sub_3241_add_2_25.INIT1 = 16'hf555;
    defparam sub_3241_add_2_25.INJECT1_0 = "NO";
    defparam sub_3241_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_23 (.A0(spi_byte_counter_31__N_760[21]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[22]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47545), .COUT(n47546));
    defparam sub_3241_add_2_23.INIT0 = 16'hf555;
    defparam sub_3241_add_2_23.INIT1 = 16'hf555;
    defparam sub_3241_add_2_23.INJECT1_0 = "NO";
    defparam sub_3241_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_21 (.A0(spi_byte_counter_31__N_760[19]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[20]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47544), .COUT(n47545));
    defparam sub_3241_add_2_21.INIT0 = 16'hf555;
    defparam sub_3241_add_2_21.INIT1 = 16'hf555;
    defparam sub_3241_add_2_21.INJECT1_0 = "NO";
    defparam sub_3241_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_19 (.A0(spi_byte_counter_31__N_760[17]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[18]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47543), .COUT(n47544));
    defparam sub_3241_add_2_19.INIT0 = 16'hf555;
    defparam sub_3241_add_2_19.INIT1 = 16'hf555;
    defparam sub_3241_add_2_19.INJECT1_0 = "NO";
    defparam sub_3241_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_17 (.A0(spi_byte_counter_31__N_760[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[16]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47542), .COUT(n47543));
    defparam sub_3241_add_2_17.INIT0 = 16'hf555;
    defparam sub_3241_add_2_17.INIT1 = 16'hf555;
    defparam sub_3241_add_2_17.INJECT1_0 = "NO";
    defparam sub_3241_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_15 (.A0(spi_byte_counter_31__N_760[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47541), .COUT(n47542));
    defparam sub_3241_add_2_15.INIT0 = 16'hf555;
    defparam sub_3241_add_2_15.INIT1 = 16'hf555;
    defparam sub_3241_add_2_15.INJECT1_0 = "NO";
    defparam sub_3241_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_13 (.A0(spi_byte_counter_31__N_760[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47540), .COUT(n47541));
    defparam sub_3241_add_2_13.INIT0 = 16'hf555;
    defparam sub_3241_add_2_13.INIT1 = 16'hf555;
    defparam sub_3241_add_2_13.INJECT1_0 = "NO";
    defparam sub_3241_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_11 (.A0(spi_byte_counter_31__N_760[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47539), .COUT(n47540));
    defparam sub_3241_add_2_11.INIT0 = 16'hf555;
    defparam sub_3241_add_2_11.INIT1 = 16'hf555;
    defparam sub_3241_add_2_11.INJECT1_0 = "NO";
    defparam sub_3241_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_9 (.A0(spi_byte_counter_31__N_760[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47538), .COUT(n47539));
    defparam sub_3241_add_2_9.INIT0 = 16'hf555;
    defparam sub_3241_add_2_9.INIT1 = 16'hf555;
    defparam sub_3241_add_2_9.INJECT1_0 = "NO";
    defparam sub_3241_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_7 (.A0(spi_byte_counter_31__N_760[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47537), .COUT(n47538));
    defparam sub_3241_add_2_7.INIT0 = 16'hf555;
    defparam sub_3241_add_2_7.INIT1 = 16'hf555;
    defparam sub_3241_add_2_7.INJECT1_0 = "NO";
    defparam sub_3241_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_5 (.A0(spi_byte_counter_31__N_760[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47536), .COUT(n47537));
    defparam sub_3241_add_2_5.INIT0 = 16'hf555;
    defparam sub_3241_add_2_5.INIT1 = 16'hf555;
    defparam sub_3241_add_2_5.INJECT1_0 = "NO";
    defparam sub_3241_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_3 (.A0(spi_byte_counter_31__N_760[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter_31__N_760[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n47535), .COUT(n47536));
    defparam sub_3241_add_2_3.INIT0 = 16'hf555;
    defparam sub_3241_add_2_3.INIT1 = 16'h0aaa;
    defparam sub_3241_add_2_3.INJECT1_0 = "NO";
    defparam sub_3241_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_3241_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter_31__N_760[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n47535));
    defparam sub_3241_add_2_1.INIT0 = 16'h0000;
    defparam sub_3241_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_3241_add_2_1.INJECT1_0 = "NO";
    defparam sub_3241_add_2_1.INJECT1_1 = "NO";
    FD1P3IX WrData_i0 (.D(WrData_23__N_691[0]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i0.GSR = "DISABLED";
    FD1P3AX SPI_CS_228 (.D(SPI_CS_N_880), .SP(sclk_c_enable_189), .CK(sclk_c), 
            .Q(CSn)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam SPI_CS_228.GSR = "DISABLED";
    FD1P3IX WrAddr_i0 (.D(WrAddr_8__N_747[0]), .SP(sclk_c_enable_1283), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(WrAddress[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i0.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i0 (.D(n1337[0]), .SP(sclk_c_enable_1315), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i0.GSR = "DISABLED";
    FD1P3IX WrEnable_i0 (.D(WrEnable_23__N_824[0]), .SP(state[0]), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(\WE[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i0.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i0 (.D(n1568[0]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i0.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i1 (.D(n1568[1]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i1.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i2 (.D(n1568[2]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i2.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i3 (.D(n1568[3]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i3.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i4 (.D(n1568[4]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i4.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i5 (.D(n1568[5]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i5.GSR = "DISABLED";
    FD1P3AY spi_byte_timeout_i6 (.D(spi_byte_timeout_31__N_595[6]), .SP(sclk_c_enable_205), 
            .CK(sclk_c), .Q(spi_byte_timeout[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i6.GSR = "DISABLED";
    FD1P3AY spi_byte_timeout_i7 (.D(spi_byte_timeout_31__N_595[7]), .SP(sclk_c_enable_205), 
            .CK(sclk_c), .Q(spi_byte_timeout[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i7.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i8 (.D(n1568[8]), .SP(sclk_c_enable_224), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(spi_byte_timeout[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i8.GSR = "DISABLED";
    FD1P3AY spi_byte_timeout_i9 (.D(spi_byte_timeout_31__N_595[9]), .SP(sclk_c_enable_205), 
            .CK(sclk_c), .Q(spi_byte_timeout[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i9.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i10 (.D(n1568[10]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i10.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i11 (.D(n1568[11]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i11.GSR = "DISABLED";
    FD1P3AY spi_byte_timeout_i12 (.D(spi_byte_timeout_31__N_595[12]), .SP(sclk_c_enable_205), 
            .CK(sclk_c), .Q(spi_byte_timeout[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i12.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i13 (.D(n1568[13]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i13.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i14 (.D(n1568[14]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i14.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i15 (.D(n1568[15]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i15.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i16 (.D(n1568[16]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i16.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i17 (.D(n1568[17]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i17.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i18 (.D(n1568[18]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i18.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i19 (.D(n1568[19]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i19.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i20 (.D(n1568[20]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i20.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i21 (.D(n1568[21]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i21.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i22 (.D(n1568[22]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i22.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i23 (.D(n1568[23]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i23.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i24 (.D(n1568[24]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i24.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i25 (.D(n1568[25]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i25.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i26 (.D(n1568[26]), .SP(sclk_c_enable_224), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_timeout[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i26.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i27 (.D(n1568[27]), .SP(sclk_c_enable_224), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_timeout[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i27.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i28 (.D(n1568[28]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i28.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i29 (.D(n1568[29]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i29.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i30 (.D(n1568[30]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i30.GSR = "DISABLED";
    FD1P3IX spi_byte_timeout_i31 (.D(n1568[31]), .SP(sclk_c_enable_224), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_timeout[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_timeout_i31.GSR = "DISABLED";
    CCU2D add_33911_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48577), 
          .S0(n14466));
    defparam add_33911_cout.INIT0 = 16'h0000;
    defparam add_33911_cout.INIT1 = 16'h0000;
    defparam add_33911_cout.INJECT1_0 = "NO";
    defparam add_33911_cout.INJECT1_1 = "NO";
    CCU2D add_33911_31 (.A0(spi_byte_timeout[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48576), .COUT(n48577));
    defparam add_33911_31.INIT0 = 16'hf555;
    defparam add_33911_31.INIT1 = 16'h5555;
    defparam add_33911_31.INJECT1_0 = "NO";
    defparam add_33911_31.INJECT1_1 = "NO";
    CCU2D add_33911_29 (.A0(spi_byte_timeout[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48575), .COUT(n48576));
    defparam add_33911_29.INIT0 = 16'hf555;
    defparam add_33911_29.INIT1 = 16'hf555;
    defparam add_33911_29.INJECT1_0 = "NO";
    defparam add_33911_29.INJECT1_1 = "NO";
    CCU2D add_33911_27 (.A0(spi_byte_timeout[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48574), .COUT(n48575));
    defparam add_33911_27.INIT0 = 16'hf555;
    defparam add_33911_27.INIT1 = 16'hf555;
    defparam add_33911_27.INJECT1_0 = "NO";
    defparam add_33911_27.INJECT1_1 = "NO";
    LUT4 mux_155_rep_1_i31_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[30]), 
         .D(n1337[30]), .Z(spi_byte_counter_31__N_760[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i31_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_143_i1_3_lut (.A(index[0]), .B(DATA_OUT[0]), .C(n14326), 
         .Z(WrAddr_8__N_747[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i1_3_lut.init = 16'hcaca;
    CCU2D add_33911_25 (.A0(spi_byte_timeout[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48573), .COUT(n48574));
    defparam add_33911_25.INIT0 = 16'hf555;
    defparam add_33911_25.INIT1 = 16'hf555;
    defparam add_33911_25.INJECT1_0 = "NO";
    defparam add_33911_25.INJECT1_1 = "NO";
    CCU2D add_33911_23 (.A0(spi_byte_timeout[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48572), .COUT(n48573));
    defparam add_33911_23.INIT0 = 16'hf555;
    defparam add_33911_23.INIT1 = 16'hf555;
    defparam add_33911_23.INJECT1_0 = "NO";
    defparam add_33911_23.INJECT1_1 = "NO";
    CCU2D add_33911_21 (.A0(spi_byte_timeout[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48571), .COUT(n48572));
    defparam add_33911_21.INIT0 = 16'hf555;
    defparam add_33911_21.INIT1 = 16'hf555;
    defparam add_33911_21.INJECT1_0 = "NO";
    defparam add_33911_21.INJECT1_1 = "NO";
    CCU2D add_33911_19 (.A0(spi_byte_timeout[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48570), .COUT(n48571));
    defparam add_33911_19.INIT0 = 16'hf555;
    defparam add_33911_19.INIT1 = 16'hf555;
    defparam add_33911_19.INJECT1_0 = "NO";
    defparam add_33911_19.INJECT1_1 = "NO";
    CCU2D add_33911_17 (.A0(spi_byte_timeout[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48569), .COUT(n48570));
    defparam add_33911_17.INIT0 = 16'hf555;
    defparam add_33911_17.INIT1 = 16'hf555;
    defparam add_33911_17.INJECT1_0 = "NO";
    defparam add_33911_17.INJECT1_1 = "NO";
    CCU2D add_33911_15 (.A0(spi_byte_timeout[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48568), .COUT(n48569));
    defparam add_33911_15.INIT0 = 16'hf555;
    defparam add_33911_15.INIT1 = 16'hf555;
    defparam add_33911_15.INJECT1_0 = "NO";
    defparam add_33911_15.INJECT1_1 = "NO";
    LUT4 mux_155_rep_1_i28_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[27]), 
         .D(n1337[27]), .Z(spi_byte_counter_31__N_760[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i28_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i29_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[28]), 
         .D(n1337[28]), .Z(spi_byte_counter_31__N_760[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i29_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i26_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[25]), 
         .D(n1337[25]), .Z(spi_byte_counter_31__N_760[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i26_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i27_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[26]), 
         .D(n1337[26]), .Z(spi_byte_counter_31__N_760[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i27_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i24_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[23]), 
         .D(n1337[23]), .Z(spi_byte_counter_31__N_760[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i24_3_lut_4_lut.init = 16'hf870;
    CCU2D add_33911_13 (.A0(spi_byte_timeout[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48567), .COUT(n48568));
    defparam add_33911_13.INIT0 = 16'hf555;
    defparam add_33911_13.INIT1 = 16'hf555;
    defparam add_33911_13.INJECT1_0 = "NO";
    defparam add_33911_13.INJECT1_1 = "NO";
    LUT4 mux_155_rep_1_i25_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[24]), 
         .D(n1337[24]), .Z(spi_byte_counter_31__N_760[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i25_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i22_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[21]), 
         .D(n1337[21]), .Z(spi_byte_counter_31__N_760[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i22_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i23_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[22]), 
         .D(n1337[22]), .Z(spi_byte_counter_31__N_760[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i23_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i20_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[19]), 
         .D(n1337[19]), .Z(spi_byte_counter_31__N_760[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i20_3_lut_4_lut.init = 16'hf870;
    CCU2D add_33911_11 (.A0(spi_byte_timeout[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48566), .COUT(n48567));
    defparam add_33911_11.INIT0 = 16'hf555;
    defparam add_33911_11.INIT1 = 16'hf555;
    defparam add_33911_11.INJECT1_0 = "NO";
    defparam add_33911_11.INJECT1_1 = "NO";
    CCU2D add_33911_9 (.A0(spi_byte_timeout[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48565), .COUT(n48566));
    defparam add_33911_9.INIT0 = 16'hf555;
    defparam add_33911_9.INIT1 = 16'hf555;
    defparam add_33911_9.INJECT1_0 = "NO";
    defparam add_33911_9.INJECT1_1 = "NO";
    LUT4 mux_206_Mux_2_i15_3_lut_4_lut (.A(index[0]), .B(index[1]), .C(index[2]), 
         .D(index[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(54[24:29])
    defparam mux_206_Mux_2_i15_3_lut_4_lut.init = 16'h9249;
    CCU2D add_33911_7 (.A0(spi_byte_timeout[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48564), .COUT(n48565));
    defparam add_33911_7.INIT0 = 16'hf555;
    defparam add_33911_7.INIT1 = 16'hf555;
    defparam add_33911_7.INJECT1_0 = "NO";
    defparam add_33911_7.INJECT1_1 = "NO";
    LUT4 mux_155_rep_1_i21_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[20]), 
         .D(n1337[20]), .Z(spi_byte_counter_31__N_760[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i21_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_206_Mux_1_i15_3_lut_4_lut (.A(index[0]), .B(index[1]), .C(index[2]), 
         .D(index[3]), .Z(n15_adj_916)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(54[24:29])
    defparam mux_206_Mux_1_i15_3_lut_4_lut.init = 16'h2492;
    LUT4 mux_206_Mux_0_i15_3_lut_4_lut (.A(index[0]), .B(index[1]), .C(index[2]), 
         .D(index[3]), .Z(n15_adj_917)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(54[24:29])
    defparam mux_206_Mux_0_i15_3_lut_4_lut.init = 16'h4924;
    LUT4 i29021_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[0]), 
         .Z(n1568[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29021_2_lut_4_lut.init = 16'h0100;
    LUT4 i29636_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[1]), 
         .Z(n1568[1])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29636_2_lut_4_lut.init = 16'h0100;
    LUT4 i29635_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[2]), 
         .Z(n1568[2])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29635_2_lut_4_lut.init = 16'h0100;
    LUT4 i29452_3_lut_4_lut (.A(index[0]), .B(index[1]), .C(index[2]), 
         .D(index[3]), .Z(n30)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(54[24:29])
    defparam i29452_3_lut_4_lut.init = 16'h0009;
    LUT4 i29634_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[3]), 
         .Z(n1568[3])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29634_2_lut_4_lut.init = 16'h0100;
    LUT4 i29633_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[4]), 
         .Z(n1568[4])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29633_2_lut_4_lut.init = 16'h0100;
    LUT4 i29632_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[5]), 
         .Z(n1568[5])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29632_2_lut_4_lut.init = 16'h0100;
    LUT4 i29631_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[8]), 
         .Z(n1568[8])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29631_2_lut_4_lut.init = 16'h0100;
    LUT4 i29630_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[10]), 
         .Z(n1568[10])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29630_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i18_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[17]), 
         .D(n1337[17]), .Z(spi_byte_counter_31__N_760[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i18_3_lut_4_lut.init = 16'hf870;
    LUT4 i29629_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[11]), 
         .Z(n1568[11])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29629_2_lut_4_lut.init = 16'h0100;
    LUT4 i29628_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[13]), 
         .Z(n1568[13])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29628_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i19_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[18]), 
         .D(n1337[18]), .Z(spi_byte_counter_31__N_760[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i19_3_lut_4_lut.init = 16'hf870;
    LUT4 i29627_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[14]), 
         .Z(n1568[14])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29627_2_lut_4_lut.init = 16'h0100;
    LUT4 i29626_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[15]), 
         .Z(n1568[15])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29626_2_lut_4_lut.init = 16'h0100;
    LUT4 i29625_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[16]), 
         .Z(n1568[16])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29625_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i16_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[15]), 
         .D(n1337[15]), .Z(spi_byte_counter_31__N_760[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i16_3_lut_4_lut.init = 16'hf870;
    LUT4 i29624_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[17]), 
         .Z(n1568[17])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29624_2_lut_4_lut.init = 16'h0100;
    CCU2D add_33911_5 (.A0(spi_byte_timeout[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48563), .COUT(n48564));
    defparam add_33911_5.INIT0 = 16'hf555;
    defparam add_33911_5.INIT1 = 16'hf555;
    defparam add_33911_5.INJECT1_0 = "NO";
    defparam add_33911_5.INJECT1_1 = "NO";
    LUT4 i29623_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[18]), 
         .Z(n1568[18])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29623_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i17_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[16]), 
         .D(n1337[16]), .Z(spi_byte_counter_31__N_760[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i17_3_lut_4_lut.init = 16'hf870;
    LUT4 i29622_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[19]), 
         .Z(n1568[19])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29622_2_lut_4_lut.init = 16'h0100;
    LUT4 i29621_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[20]), 
         .Z(n1568[20])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29621_2_lut_4_lut.init = 16'h0100;
    LUT4 i29620_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[21]), 
         .Z(n1568[21])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29620_2_lut_4_lut.init = 16'h0100;
    LUT4 i29619_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[22]), 
         .Z(n1568[22])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29619_2_lut_4_lut.init = 16'h0100;
    LUT4 i29618_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[23]), 
         .Z(n1568[23])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29618_2_lut_4_lut.init = 16'h0100;
    LUT4 i29617_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[24]), 
         .Z(n1568[24])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29617_2_lut_4_lut.init = 16'h0100;
    LUT4 i29616_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[25]), 
         .Z(n1568[25])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29616_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i14_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[13]), 
         .D(n1337[13]), .Z(spi_byte_counter_31__N_760[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i14_3_lut_4_lut.init = 16'hf870;
    LUT4 i29615_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[26]), 
         .Z(n1568[26])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29615_2_lut_4_lut.init = 16'h0100;
    LUT4 i29614_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[27]), 
         .Z(n1568[27])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29614_2_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut (.A(sclk_c_enable_224), .B(n55545), .Z(sclk_c_enable_205)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i29613_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[28]), 
         .Z(n1568[28])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29613_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i15_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[14]), 
         .D(n1337[14]), .Z(spi_byte_counter_31__N_760[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i15_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i12_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[11]), 
         .D(n1337[11]), .Z(spi_byte_counter_31__N_760[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i12_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i13_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[12]), 
         .D(n1337[12]), .Z(spi_byte_counter_31__N_760[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i13_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_3_lut (.A(n98), .B(n44072), .C(n869[6]), .Z(spi_byte_timeout_31__N_595[6])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i29612_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[29]), 
         .Z(n1568[29])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29612_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i10_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[9]), 
         .D(n1337[9]), .Z(spi_byte_counter_31__N_760[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i10_3_lut_4_lut.init = 16'hf870;
    LUT4 i29611_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[30]), 
         .Z(n1568[30])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29611_2_lut_4_lut.init = 16'h0100;
    LUT4 mux_155_rep_1_i11_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[10]), 
         .D(n1337[10]), .Z(spi_byte_counter_31__N_760[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i11_3_lut_4_lut.init = 16'hf870;
    LUT4 i29610_2_lut_4_lut (.A(n14501), .B(RX_RDY), .C(n14466), .D(n869[31]), 
         .Z(n1568[31])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29610_2_lut_4_lut.init = 16'h0100;
    LUT4 i31971_3_lut (.A(n54553), .B(n55544), .C(n55545), .Z(n44072)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i31971_3_lut.init = 16'h3a3a;
    LUT4 mux_155_rep_1_i8_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[7]), 
         .D(n1337[7]), .Z(spi_byte_counter_31__N_760[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i8_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_3_lut_adj_842 (.A(n98), .B(n44072), .C(n869[7]), .Z(spi_byte_timeout_31__N_595[7])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_adj_842.init = 16'hecec;
    LUT4 mux_155_rep_1_i9_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[8]), 
         .D(n1337[8]), .Z(spi_byte_counter_31__N_760[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i9_3_lut_4_lut.init = 16'hf870;
    LUT4 i38536_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8), 
         .Z(WrEnable_23__N_824[19])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38536_2_lut_2_lut_4_lut.init = 16'h0040;
    LUT4 i38524_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_918), 
         .Z(WrEnable_23__N_824[15])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38524_2_lut_2_lut_4_lut.init = 16'h0040;
    LUT4 mux_155_rep_1_i6_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[5]), 
         .D(n1337[5]), .Z(spi_byte_counter_31__N_760[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i6_3_lut_4_lut.init = 16'hf870;
    LUT4 i38512_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_919), 
         .Z(WrEnable_23__N_824[11])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38512_2_lut_2_lut_4_lut.init = 16'h0040;
    LUT4 i38500_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_920), 
         .Z(WrEnable_23__N_824[7])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38500_2_lut_2_lut_4_lut.init = 16'h0040;
    LUT4 mux_155_rep_1_i7_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[6]), 
         .D(n1337[6]), .Z(spi_byte_counter_31__N_760[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i7_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_3_lut_adj_843 (.A(n98), .B(n44072), .C(n869[9]), .Z(spi_byte_timeout_31__N_595[9])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_adj_843.init = 16'hecec;
    LUT4 i38488_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_921), 
         .Z(WrEnable_23__N_824[3])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38488_2_lut_2_lut_4_lut.init = 16'h0040;
    LUT4 mux_155_rep_1_i4_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[3]), 
         .D(n1337[3]), .Z(spi_byte_counter_31__N_760[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i4_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_155_rep_1_i5_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[4]), 
         .D(n1337[4]), .Z(spi_byte_counter_31__N_760[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i5_3_lut_4_lut.init = 16'hf870;
    CCU2D add_33911_3 (.A0(spi_byte_timeout[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48562), .COUT(n48563));
    defparam add_33911_3.INIT0 = 16'hf555;
    defparam add_33911_3.INIT1 = 16'hf555;
    defparam add_33911_3.INJECT1_0 = "NO";
    defparam add_33911_3.INJECT1_1 = "NO";
    LUT4 i38533_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8), 
         .Z(WrEnable_23__N_824[18])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i38533_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 mux_155_rep_1_i2_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[1]), 
         .D(n1337[1]), .Z(spi_byte_counter_31__N_760[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i2_3_lut_4_lut.init = 16'hf870;
    LUT4 i38521_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_918), 
         .Z(WrEnable_23__N_824[14])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i38521_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 mux_155_rep_1_i3_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[2]), 
         .D(n1337[2]), .Z(spi_byte_counter_31__N_760[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i3_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_3_lut_adj_844 (.A(n98), .B(n44072), .C(n869[12]), .Z(spi_byte_timeout_31__N_595[12])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_adj_844.init = 16'hecec;
    LUT4 i38509_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_919), 
         .Z(WrEnable_23__N_824[10])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i38509_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 i38497_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_920), 
         .Z(WrEnable_23__N_824[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i38497_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 i38485_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_921), 
         .Z(WrEnable_23__N_824[2])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i38485_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 i38530_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8), 
         .Z(WrEnable_23__N_824[17])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i38530_2_lut_2_lut_4_lut.init = 16'h0004;
    LUT4 i38518_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_918), 
         .Z(WrEnable_23__N_824[13])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i38518_2_lut_2_lut_4_lut.init = 16'h0004;
    LUT4 mux_155_rep_1_i1_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[0]), 
         .D(n1337[0]), .Z(spi_byte_counter_31__N_760[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i1_3_lut_4_lut.init = 16'hf870;
    LUT4 i38568_2_lut_3_lut (.A(n14326), .B(n54553), .C(n55544), .Z(sclk_c_enable_1315)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i38568_2_lut_3_lut.init = 16'h0808;
    LUT4 i38506_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_919), 
         .Z(WrEnable_23__N_824[9])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i38506_2_lut_2_lut_4_lut.init = 16'h0004;
    LUT4 i38494_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_920), 
         .Z(WrEnable_23__N_824[5])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i38494_2_lut_2_lut_4_lut.init = 16'h0004;
    LUT4 i38482_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_921), 
         .Z(WrEnable_23__N_824[1])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i38482_2_lut_2_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut (.A(fb[3]), .B(fb[4]), .C(fb[2]), .Z(n8)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i38539_3_lut_4_lut (.A(fb[3]), .B(fb[4]), .C(n54678), .D(fb[2]), 
         .Z(WrEnable_23__N_824[20])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i38539_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_adj_845 (.A(fb[4]), .B(fb[2]), .C(fb[3]), .Z(n8_adj_920)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i1_2_lut_3_lut_adj_845.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_846 (.A(fb[4]), .B(fb[2]), .C(fb[3]), .Z(n8_adj_918)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i1_2_lut_3_lut_adj_846.init = 16'hbfbf;
    LUT4 i2_4_lut_then_4_lut (.A(n14326), .B(n51598), .C(n14361), .D(n55544), 
         .Z(n55003)) /* synthesis lut_function=(!((B ((D)+!C)+!B (D))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i2_4_lut_then_4_lut.init = 16'h00a2;
    LUT4 i2_4_lut_else_4_lut (.A(n14326), .B(n14501), .C(n55544), .Z(n55002)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i2_4_lut_else_4_lut.init = 16'h0202;
    CCU2D add_33911_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(spi_byte_timeout[0]), .B1(spi_byte_timeout[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48562));
    defparam add_33911_1.INIT0 = 16'hF000;
    defparam add_33911_1.INIT1 = 16'ha666;
    defparam add_33911_1.INJECT1_0 = "NO";
    defparam add_33911_1.INJECT1_1 = "NO";
    FD1P3AX delay_counter_i31 (.D(delay_counter_31__N_531[31]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i31.GSR = "DISABLED";
    FD1P3AX delay_counter_i30 (.D(delay_counter_31__N_531[30]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i30.GSR = "DISABLED";
    FD1P3AX delay_counter_i29 (.D(delay_counter_31__N_531[29]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i29.GSR = "DISABLED";
    FD1P3AX delay_counter_i28 (.D(delay_counter_31__N_531[28]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i28.GSR = "DISABLED";
    FD1P3AX delay_counter_i27 (.D(delay_counter_31__N_531[27]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i27.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(RX_RDY), .B(n54680), .C(n55545), .D(n14501), 
         .Z(n98)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i2_3_lut_4_lut.init = 16'h000d;
    FD1P3AX delay_counter_i26 (.D(delay_counter_31__N_531[26]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i26.GSR = "DISABLED";
    FD1P3AX delay_counter_i25 (.D(delay_counter_31__N_531[25]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i25.GSR = "DISABLED";
    FD1P3AX delay_counter_i24 (.D(delay_counter_31__N_531[24]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i24.GSR = "DISABLED";
    FD1P3AX delay_counter_i23 (.D(delay_counter_31__N_531[23]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i23.GSR = "DISABLED";
    FD1P3AX delay_counter_i22 (.D(delay_counter_31__N_531[22]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i22.GSR = "DISABLED";
    FD1P3AX delay_counter_i21 (.D(delay_counter_31__N_531[21]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i21.GSR = "DISABLED";
    FD1P3AX delay_counter_i20 (.D(delay_counter_31__N_531[20]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i20.GSR = "DISABLED";
    FD1P3AX delay_counter_i19 (.D(delay_counter_31__N_531[19]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i19.GSR = "DISABLED";
    FD1P3AX delay_counter_i18 (.D(delay_counter_31__N_531[18]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i18.GSR = "DISABLED";
    FD1P3AX delay_counter_i17 (.D(delay_counter_31__N_531[17]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i17.GSR = "DISABLED";
    FD1P3AX delay_counter_i16 (.D(delay_counter_31__N_531[16]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i16.GSR = "DISABLED";
    FD1P3AX delay_counter_i15 (.D(delay_counter_31__N_531[15]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i15.GSR = "DISABLED";
    FD1P3AX delay_counter_i14 (.D(delay_counter_31__N_531[14]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i14.GSR = "DISABLED";
    FD1P3AX delay_counter_i13 (.D(delay_counter_31__N_531[13]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i13.GSR = "DISABLED";
    FD1P3AX delay_counter_i12 (.D(delay_counter_31__N_531[12]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i12.GSR = "DISABLED";
    FD1P3AX delay_counter_i11 (.D(delay_counter_31__N_531[11]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i11.GSR = "DISABLED";
    FD1P3AX delay_counter_i10 (.D(delay_counter_31__N_531[10]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i10.GSR = "DISABLED";
    FD1P3AX delay_counter_i9 (.D(delay_counter_31__N_531[9]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i8 (.D(delay_counter_31__N_531[8]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i7 (.D(delay_counter_31__N_531[7]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i6 (.D(delay_counter_31__N_531[6]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i6.GSR = "DISABLED";
    FD1P3AX delay_counter_i5 (.D(delay_counter_31__N_531[5]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i5.GSR = "DISABLED";
    FD1P3AX delay_counter_i4 (.D(delay_counter_31__N_531[4]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i4.GSR = "DISABLED";
    FD1P3AX delay_counter_i3 (.D(delay_counter_31__N_531[3]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i3.GSR = "DISABLED";
    FD1P3IX delay_counter_i2 (.D(n1), .SP(sclk_c_enable_1027), .CD(n36657), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i2.GSR = "DISABLED";
    FD1P3AX delay_counter_i1 (.D(delay_counter_31__N_531[1]), .SP(sclk_c_enable_1027), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i1.GSR = "DISABLED";
    FD1P3IX index_i31 (.D(index_31__N_848[31]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i31.GSR = "DISABLED";
    FD1P3IX index_i30 (.D(index_31__N_848[30]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i30.GSR = "DISABLED";
    FD1P3IX index_i29 (.D(index_31__N_848[29]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i29.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_675 (.A(n14571), .B(fb[0]), .C(fb[1]), .Z(n54678)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_675.init = 16'hfefe;
    LUT4 i38515_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_918), 
         .Z(WrEnable_23__N_824[12])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38515_2_lut_2_lut_4_lut.init = 16'h0001;
    LUT4 i38527_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8), 
         .Z(WrEnable_23__N_824[16])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38527_2_lut_2_lut_4_lut.init = 16'h0001;
    FD1P3IX index_i28 (.D(index_31__N_848[28]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i28.GSR = "DISABLED";
    LUT4 i38503_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_919), 
         .Z(WrEnable_23__N_824[8])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38503_2_lut_2_lut_4_lut.init = 16'h0001;
    FD1P3IX index_i27 (.D(index_31__N_848[27]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i27.GSR = "DISABLED";
    FD1P3IX index_i26 (.D(index_31__N_848[26]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i26.GSR = "DISABLED";
    FD1P3IX index_i25 (.D(index_31__N_848[25]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i25.GSR = "DISABLED";
    FD1P3IX index_i24 (.D(index_31__N_848[24]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i24.GSR = "DISABLED";
    LUT4 i38491_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_920), 
         .Z(WrEnable_23__N_824[4])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38491_2_lut_2_lut_4_lut.init = 16'h0001;
    LUT4 i38456_2_lut_2_lut_4_lut (.A(n14571), .B(fb[0]), .C(fb[1]), .D(n8_adj_921), 
         .Z(WrEnable_23__N_824[0])) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38456_2_lut_2_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_rep_676 (.A(RX_RDY), .B(n14361), .Z(n54679)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_2_lut_rep_676.init = 16'h8888;
    LUT4 i1_2_lut_rep_619_3_lut (.A(RX_RDY), .B(n14361), .C(n14396), .Z(n54622)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_2_lut_rep_619_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(RX_RDY), .B(n14361), .C(n14431), .D(n14396), 
         .Z(n131)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3IX index_i23 (.D(index_31__N_848[23]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0 (.D(n1_adj_922), .SP(sclk_c_enable_1027), .CD(n36657), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam delay_counter_i0.GSR = "DISABLED";
    FD1P3IX index_i0 (.D(index_31__N_848[0]), .SP(sclk_c_enable_1028), .CD(n36657), 
            .CK(sclk_c), .Q(index[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i0.GSR = "DISABLED";
    FD1P3IX index_i22 (.D(index_31__N_848[22]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i22.GSR = "DISABLED";
    FD1P3IX index_i21 (.D(index_31__N_848[21]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i21.GSR = "DISABLED";
    FD1P3IX index_i20 (.D(index_31__N_848[20]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i20.GSR = "DISABLED";
    FD1P3IX index_i19 (.D(index_31__N_848[19]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i19.GSR = "DISABLED";
    FD1P3IX index_i18 (.D(index_31__N_848[18]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i18.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_625_4_lut (.A(RX_RDY), .B(n14361), .C(n14326), .D(n14396), 
         .Z(n54628)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_3_lut_rep_625_4_lut.init = 16'h0f8f;
    LUT4 i1_2_lut_rep_677 (.A(n14361), .B(n51598), .Z(n54680)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_677.init = 16'hbbbb;
    LUT4 i29041_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[17]), 
         .D(RX_RDY), .Z(n1337[17])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29041_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29025_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[1]), 
         .D(RX_RDY), .Z(n1337[1])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29025_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29043_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[19]), 
         .D(RX_RDY), .Z(n1337[19])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29043_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29044_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[20]), 
         .D(RX_RDY), .Z(n1337[20])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29044_2_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3IX state_i0 (.D(n1_adj_923), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3IX fb_i0 (.D(fb_31__N_715[0]), .SP(sclk_c_enable_1111), .CD(n36653), 
            .CK(sclk_c), .Q(fb[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam fb_i0.GSR = "DISABLED";
    FD1P3IX index_i17 (.D(index_31__N_848[17]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i17.GSR = "DISABLED";
    LUT4 i29053_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[29]), 
         .D(RX_RDY), .Z(n1337[29])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29053_2_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3IX index_i16 (.D(index_31__N_848[16]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i16.GSR = "DISABLED";
    FD1P3IX index_i15 (.D(index_31__N_848[15]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i15.GSR = "DISABLED";
    FD1P3IX index_i14 (.D(index_31__N_848[14]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i14.GSR = "DISABLED";
    FD1P3IX index_i13 (.D(index_31__N_848[13]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i13.GSR = "DISABLED";
    LUT4 i29046_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[22]), 
         .D(RX_RDY), .Z(n1337[22])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29046_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29045_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[21]), 
         .D(RX_RDY), .Z(n1337[21])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29045_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29047_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[23]), 
         .D(RX_RDY), .Z(n1337[23])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29047_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29048_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[24]), 
         .D(RX_RDY), .Z(n1337[24])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29048_2_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3IX index_i12 (.D(index_31__N_848[12]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i12.GSR = "DISABLED";
    FD1P3IX index_i11 (.D(index_31__N_848[11]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i11.GSR = "DISABLED";
    FD1P3IX index_i10 (.D(index_31__N_848[10]), .SP(sclk_c_enable_1092), 
            .CD(n36657), .CK(sclk_c), .Q(index[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i10.GSR = "DISABLED";
    FD1P3IX index_i9 (.D(index_31__N_848[9]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i9.GSR = "DISABLED";
    FD1P3IX index_i8 (.D(index_31__N_848[8]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i8.GSR = "DISABLED";
    FD1P3IX index_i7 (.D(index_31__N_848[7]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i7.GSR = "DISABLED";
    FD1P3IX index_i6 (.D(index_31__N_848[6]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i6.GSR = "DISABLED";
    FD1P3IX index_i5 (.D(index_31__N_848[5]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i5.GSR = "DISABLED";
    LUT4 i29050_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[26]), 
         .D(RX_RDY), .Z(n1337[26])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29050_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29049_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[25]), 
         .D(RX_RDY), .Z(n1337[25])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29049_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29052_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[28]), 
         .D(RX_RDY), .Z(n1337[28])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29052_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29051_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[27]), 
         .D(RX_RDY), .Z(n1337[27])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29051_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29054_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[30]), 
         .D(RX_RDY), .Z(n1337[30])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29054_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29055_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[31]), 
         .D(RX_RDY), .Z(n1337[31])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29055_2_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3IX index_i4 (.D(index_31__N_848[4]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i4.GSR = "DISABLED";
    FD1P3IX index_i3 (.D(index_31__N_848[3]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i3.GSR = "DISABLED";
    FD1P3IX index_i2 (.D(index_31__N_848[2]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i2.GSR = "DISABLED";
    FD1P3IX index_i1 (.D(index_31__N_848[1]), .SP(sclk_c_enable_1092), .CD(n36657), 
            .CK(sclk_c), .Q(index[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam index_i1.GSR = "DISABLED";
    FD1P3IX state_i1 (.D(state[0]), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3IX fb_i4 (.D(fb_31__N_715[4]), .SP(sclk_c_enable_1111), .CD(n36653), 
            .CK(sclk_c), .Q(fb[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam fb_i4.GSR = "DISABLED";
    LUT4 i28670_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[0]), 
         .D(RX_RDY), .Z(n1337[0])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i28670_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29042_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[18]), 
         .D(RX_RDY), .Z(n1337[18])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29042_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29040_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[16]), 
         .D(RX_RDY), .Z(n1337[16])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29040_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29039_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[15]), 
         .D(RX_RDY), .Z(n1337[15])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29039_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29037_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[13]), 
         .D(RX_RDY), .Z(n1337[13])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29037_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29038_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[14]), 
         .D(RX_RDY), .Z(n1337[14])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29038_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29035_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[11]), 
         .D(RX_RDY), .Z(n1337[11])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29035_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29036_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[12]), 
         .D(RX_RDY), .Z(n1337[12])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29036_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29034_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[10]), 
         .D(RX_RDY), .Z(n1337[10])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29034_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29033_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[9]), 
         .D(RX_RDY), .Z(n1337[9])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29033_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29031_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[7]), 
         .D(RX_RDY), .Z(n1337[7])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29031_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29032_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[8]), 
         .D(RX_RDY), .Z(n1337[8])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29032_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29030_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[6]), 
         .D(RX_RDY), .Z(n1337[6])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29030_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29029_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[5]), 
         .D(RX_RDY), .Z(n1337[5])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29029_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29027_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[3]), 
         .D(RX_RDY), .Z(n1337[3])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29027_2_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3IX fb_i3 (.D(fb_31__N_715[3]), .SP(sclk_c_enable_1111), .CD(n36653), 
            .CK(sclk_c), .Q(fb[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam fb_i3.GSR = "DISABLED";
    FD1P3IX fb_i2 (.D(fb_31__N_715[2]), .SP(sclk_c_enable_1111), .CD(n36653), 
            .CK(sclk_c), .Q(fb[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam fb_i2.GSR = "DISABLED";
    FD1P3IX fb_i1 (.D(fb_31__N_715[1]), .SP(sclk_c_enable_1111), .CD(n36653), 
            .CK(sclk_c), .Q(fb[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam fb_i1.GSR = "DISABLED";
    LUT4 i29028_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[4]), 
         .D(RX_RDY), .Z(n1337[4])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29028_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i29026_2_lut_3_lut_4_lut (.A(n14361), .B(n51598), .C(n830[2]), 
         .D(RX_RDY), .Z(n1337[2])) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i29026_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i1_3_lut_4_lut (.A(n54742), .B(n14326), .C(n51592), .D(spi_byte_counter[0]), 
         .Z(sclk_c_enable_1260)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_4_lut.init = 16'hf111;
    LUT4 i1_3_lut_4_lut_adj_847 (.A(n54742), .B(n14326), .C(n51592), .D(spi_byte_counter[0]), 
         .Z(sclk_c_enable_1268)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_4_lut_adj_847.init = 16'h11f1;
    FD1P3IX WrData_i1 (.D(WrData_23__N_691[1]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i1.GSR = "DISABLED";
    FD1P3IX WrData_i2 (.D(WrData_23__N_691[2]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i2.GSR = "DISABLED";
    FD1P3IX WrData_i3 (.D(WrData_23__N_691[3]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i3.GSR = "DISABLED";
    FD1P3IX WrData_i4 (.D(WrData_23__N_691[4]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i4.GSR = "DISABLED";
    FD1P3IX WrData_i5 (.D(WrData_23__N_691[5]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i5.GSR = "DISABLED";
    FD1P3IX WrData_i6 (.D(WrData_23__N_691[6]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i6.GSR = "DISABLED";
    FD1P3IX WrData_i7 (.D(WrData_23__N_691[7]), .SP(sclk_c_enable_1260), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i7.GSR = "DISABLED";
    FD1P3IX WrData_i8 (.D(WrData_23__N_691[8]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i8.GSR = "DISABLED";
    FD1P3IX WrData_i9 (.D(WrData_23__N_691[9]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[9])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i9.GSR = "DISABLED";
    FD1P3IX WrData_i10 (.D(WrData_23__N_691[10]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[10])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i10.GSR = "DISABLED";
    FD1P3IX WrData_i11 (.D(WrData_23__N_691[11]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[11])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i11.GSR = "DISABLED";
    FD1P3IX WrData_i12 (.D(WrData_23__N_691[12]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[12])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i12.GSR = "DISABLED";
    FD1P3IX WrData_i13 (.D(WrData_23__N_691[13]), .SP(sclk_c_enable_1268), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(Data[13])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i13.GSR = "DISABLED";
    FD1P3IX WrData_i14 (.D(WrData_23__N_691[14]), .SP(sclk_c_enable_1268), 
            .CD(n55547), .CK(sclk_c), .Q(Data[14])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i14.GSR = "DISABLED";
    FD1P3IX WrData_i15 (.D(WrData_23__N_691[15]), .SP(sclk_c_enable_1268), 
            .CD(n55547), .CK(sclk_c), .Q(Data[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i15.GSR = "DISABLED";
    FD1P3IX WrData_i16 (.D(WrData_23__N_691[16]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[16])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i16.GSR = "DISABLED";
    FD1P3IX WrData_i17 (.D(WrData_23__N_691[17]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[17])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i17.GSR = "DISABLED";
    FD1P3IX WrData_i18 (.D(WrData_23__N_691[18]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[18])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i18.GSR = "DISABLED";
    FD1P3IX WrData_i19 (.D(WrData_23__N_691[19]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[19])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i19.GSR = "DISABLED";
    FD1P3IX WrData_i20 (.D(WrData_23__N_691[20]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[20])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i20.GSR = "DISABLED";
    FD1P3IX WrData_i21 (.D(WrData_23__N_691[21]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[21])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i21.GSR = "DISABLED";
    FD1P3IX WrData_i22 (.D(WrData_23__N_691[22]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[22])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i22.GSR = "DISABLED";
    FD1P3IX WrData_i23 (.D(WrData_23__N_691[23]), .SP(sclk_c_enable_1276), 
            .CD(n55547), .CK(sclk_c), .Q(Data[23])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrData_i23.GSR = "DISABLED";
    FD1P3IX WrAddr_i1 (.D(WrAddr_8__N_747[1]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i1.GSR = "DISABLED";
    FD1P3IX WrAddr_i2 (.D(WrAddr_8__N_747[2]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i2.GSR = "DISABLED";
    FD1P3IX WrAddr_i3 (.D(WrAddr_8__N_747[3]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i3.GSR = "DISABLED";
    FD1P3IX WrAddr_i4 (.D(WrAddr_8__N_747[4]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i4.GSR = "DISABLED";
    FD1P3IX WrAddr_i5 (.D(WrAddr_8__N_747[5]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i5.GSR = "DISABLED";
    FD1P3IX WrAddr_i6 (.D(WrAddr_8__N_747[6]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i6.GSR = "DISABLED";
    FD1P3IX WrAddr_i7 (.D(WrAddr_8__N_747[7]), .SP(sclk_c_enable_1283), 
            .CD(n55547), .CK(sclk_c), .Q(WrAddress[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i7.GSR = "DISABLED";
    FD1P3IX WrAddr_i8 (.D(WrAddr_8__N_747[8]), .SP(sclk_c_enable_1284), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(WrAddress[8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrAddr_i8.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i1 (.D(n1337[1]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i1.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i2 (.D(n1337[2]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i2.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i3 (.D(n1337[3]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i3.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i4 (.D(n1337[4]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i4.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i5 (.D(n1337[5]), .SP(sclk_c_enable_1315), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i5.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i6 (.D(n1337[6]), .SP(sclk_c_enable_1315), 
            .CD(sclk_c_enable_1028), .CK(sclk_c), .Q(spi_byte_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i6.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i7 (.D(n1337[7]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i7.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i8 (.D(n1337[8]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i8.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i9 (.D(n1337[9]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i9.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i10 (.D(n1337[10]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i10.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i11 (.D(n1337[11]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i11.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i12 (.D(n1337[12]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i12.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i13 (.D(n1337[13]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i13.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i14 (.D(n1337[14]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i14.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i15 (.D(n1337[15]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i15.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i16 (.D(n1337[16]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i16.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i17 (.D(n1337[17]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i17.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i18 (.D(n1337[18]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i18.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i19 (.D(n1337[19]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i19.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i20 (.D(n1337[20]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i20.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i21 (.D(n1337[21]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i21.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i22 (.D(n1337[22]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i22.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i23 (.D(n1337[23]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i23.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i24 (.D(n1337[24]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i24.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i25 (.D(n1337[25]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i25.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i26 (.D(n1337[26]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i26.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i27 (.D(n1337[27]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i27.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i28 (.D(n1337[28]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i28.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i29 (.D(n1337[29]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i29.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i30 (.D(n1337[30]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i30.GSR = "DISABLED";
    FD1P3IX spi_byte_counter_i31 (.D(n1337[31]), .SP(sclk_c_enable_1315), 
            .CD(n55547), .CK(sclk_c), .Q(spi_byte_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam spi_byte_counter_i31.GSR = "DISABLED";
    FD1P3IX WrEnable_i1 (.D(WrEnable_23__N_824[1]), .SP(state[0]), .CD(n55547), 
            .CK(sclk_c), .Q(\WE[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i1.GSR = "DISABLED";
    FD1P3IX WrEnable_i2 (.D(WrEnable_23__N_824[2]), .SP(state[0]), .CD(n55547), 
            .CK(sclk_c), .Q(\WE[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i2.GSR = "DISABLED";
    FD1P3IX WrEnable_i3 (.D(WrEnable_23__N_824[3]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i3.GSR = "DISABLED";
    FD1P3IX WrEnable_i4 (.D(WrEnable_23__N_824[4]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i4.GSR = "DISABLED";
    FD1P3IX WrEnable_i5 (.D(WrEnable_23__N_824[5]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i5.GSR = "DISABLED";
    FD1P3IX WrEnable_i6 (.D(WrEnable_23__N_824[6]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i6.GSR = "DISABLED";
    FD1P3IX WrEnable_i7 (.D(WrEnable_23__N_824[7]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i7.GSR = "DISABLED";
    FD1P3IX WrEnable_i8 (.D(WrEnable_23__N_824[8]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i8.GSR = "DISABLED";
    FD1P3IX WrEnable_i9 (.D(WrEnable_23__N_824[9]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[9] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i9.GSR = "DISABLED";
    FD1P3IX WrEnable_i10 (.D(WrEnable_23__N_824[10]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i10.GSR = "DISABLED";
    FD1P3IX WrEnable_i11 (.D(WrEnable_23__N_824[11]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i11.GSR = "DISABLED";
    FD1P3IX WrEnable_i12 (.D(WrEnable_23__N_824[12]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i12.GSR = "DISABLED";
    FD1P3IX WrEnable_i13 (.D(WrEnable_23__N_824[13]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[13] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i13.GSR = "DISABLED";
    FD1P3IX WrEnable_i14 (.D(WrEnable_23__N_824[14]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[14] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i14.GSR = "DISABLED";
    FD1P3IX WrEnable_i15 (.D(WrEnable_23__N_824[15]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[15] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i15.GSR = "DISABLED";
    FD1P3IX WrEnable_i16 (.D(WrEnable_23__N_824[16]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[16] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i16.GSR = "DISABLED";
    FD1P3IX WrEnable_i17 (.D(WrEnable_23__N_824[17]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[17] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i17.GSR = "DISABLED";
    FD1P3IX WrEnable_i18 (.D(WrEnable_23__N_824[18]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[18] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i18.GSR = "DISABLED";
    FD1P3IX WrEnable_i19 (.D(WrEnable_23__N_824[19]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[19] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i19.GSR = "DISABLED";
    FD1P3IX WrEnable_i20 (.D(WrEnable_23__N_824[20]), .SP(state[0]), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(\WE[20] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam WrEnable_i20.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_848 (.A(fb[4]), .B(fb[2]), .C(fb[3]), .Z(n8_adj_921)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i1_2_lut_3_lut_adj_848.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_849 (.A(fb[4]), .B(fb[2]), .C(fb[3]), .Z(n8_adj_919)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(96[14:16])
    defparam i1_2_lut_3_lut_adj_849.init = 16'hefef;
    LUT4 mux_155_rep_1_i30_3_lut_4_lut (.A(n14326), .B(n54553), .C(spi_byte_counter[29]), 
         .D(n1337[29]), .Z(spi_byte_counter_31__N_760[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_155_rep_1_i30_3_lut_4_lut.init = 16'hf870;
    LUT4 i4_4_lut (.A(DATA_OUT[4]), .B(n52919), .C(DATA_OUT[6]), .D(n6), 
         .Z(n51598)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i4_4_lut.init = 16'hfffb;
    LUT4 i37713_4_lut (.A(DATA_OUT[0]), .B(DATA_OUT[2]), .C(DATA_OUT[1]), 
         .D(DATA_OUT[3]), .Z(n52919)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i37713_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_850 (.A(DATA_OUT[5]), .B(DATA_OUT[7]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_850.init = 16'heeee;
    LUT4 i1_3_lut_rep_550_4_lut_then_3_lut (.A(n51598), .B(n14361), .C(RX_RDY), 
         .Z(n54881)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_3_lut_rep_550_4_lut_then_3_lut.init = 16'hd0d0;
    LUT4 i1_3_lut_rep_550_4_lut_else_3_lut (.A(n51598), .B(n14361), .C(n14466), 
         .D(RX_RDY), .Z(n54880)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C+(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(113[12:18])
    defparam i1_3_lut_rep_550_4_lut_else_3_lut.init = 16'hddf0;
    LUT4 mux_129_i2_3_lut (.A(n2[7]), .B(DATA_OUT[1]), .C(n14326), .Z(WrData_23__N_691[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i2_3_lut.init = 16'hcaca;
    LUT4 mux_129_i3_3_lut (.A(n2[7]), .B(DATA_OUT[2]), .C(n14326), .Z(WrData_23__N_691[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i3_3_lut.init = 16'hcaca;
    LUT4 mux_129_i4_3_lut (.A(n2[7]), .B(DATA_OUT[3]), .C(n14326), .Z(WrData_23__N_691[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i4_3_lut.init = 16'hcaca;
    LUT4 mux_129_i5_3_lut (.A(n2[7]), .B(DATA_OUT[4]), .C(n14326), .Z(WrData_23__N_691[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i5_3_lut.init = 16'hcaca;
    LUT4 mux_129_i6_3_lut (.A(n2[7]), .B(DATA_OUT[5]), .C(n14326), .Z(WrData_23__N_691[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i6_3_lut.init = 16'hcaca;
    LUT4 mux_129_i7_3_lut (.A(n2[7]), .B(DATA_OUT[6]), .C(n14326), .Z(WrData_23__N_691[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i7_3_lut.init = 16'hcaca;
    LUT4 mux_129_i8_3_lut (.A(n2[7]), .B(DATA_OUT[7]), .C(n14326), .Z(WrData_23__N_691[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i8_3_lut.init = 16'hcaca;
    LUT4 mux_129_i9_3_lut (.A(n2[15]), .B(DATA_OUT[0]), .C(n14326), .Z(WrData_23__N_691[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i9_3_lut.init = 16'hcaca;
    LUT4 mux_129_i10_3_lut (.A(n2[15]), .B(DATA_OUT[1]), .C(n14326), .Z(WrData_23__N_691[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i10_3_lut.init = 16'hcaca;
    LUT4 mux_129_i11_3_lut (.A(n2[15]), .B(DATA_OUT[2]), .C(n14326), .Z(WrData_23__N_691[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i11_3_lut.init = 16'hcaca;
    LUT4 mux_129_i12_3_lut (.A(n2[15]), .B(DATA_OUT[3]), .C(n14326), .Z(WrData_23__N_691[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i12_3_lut.init = 16'hcaca;
    LUT4 mux_129_i13_3_lut (.A(n2[15]), .B(DATA_OUT[4]), .C(n14326), .Z(WrData_23__N_691[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i13_3_lut.init = 16'hcaca;
    LUT4 mux_129_i14_3_lut (.A(n2[15]), .B(DATA_OUT[5]), .C(n14326), .Z(WrData_23__N_691[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i14_3_lut.init = 16'hcaca;
    LUT4 mux_129_i15_3_lut (.A(n2[15]), .B(DATA_OUT[6]), .C(n14326), .Z(WrData_23__N_691[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_737 (.A(n55544), .B(n55545), .Z(sclk_c_enable_1027)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_737.init = 16'hbbbb;
    LUT4 mux_129_i16_3_lut (.A(n2[15]), .B(DATA_OUT[7]), .C(n14326), .Z(WrData_23__N_691[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i16_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_738 (.A(n55545), .B(n55544), .Z(n54741)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_2_lut_rep_738.init = 16'hbbbb;
    LUT4 i1_3_lut_4_lut_adj_851 (.A(n55545), .B(n55544), .C(n49273), .D(n14326), 
         .Z(sclk_c_enable_1276)) /* synthesis lut_function=(A (C+!(D))+!A !(B+!(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_3_lut_4_lut_adj_851.init = 16'hb0bb;
    LUT4 i2_4_lut_rep_563_4_lut_3_lut (.A(n55545), .B(n55544), .C(n54628), 
         .Z(sclk_c_enable_1111)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i2_4_lut_rep_563_4_lut_3_lut.init = 16'h9898;
    LUT4 i1_2_lut_3_lut_2_lut (.A(n55545), .B(n55544), .Z(sclk_c_enable_189)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_2_lut_3_lut_2_lut.init = 16'h9999;
    LUT4 i24443_2_lut_3_lut_3_lut_2_lut (.A(n55545), .B(n55544), .Z(n36653)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i24443_2_lut_3_lut_3_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_739 (.A(n55544), .B(n55545), .Z(n54742)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_rep_739.init = 16'h2222;
    LUT4 i1_2_lut_rep_678_3_lut (.A(n55544), .B(n55545), .C(n14326), .Z(n54681)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_rep_678_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut_adj_852 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[31]), 
         .Z(delay_counter_31__N_531[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_852.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_853 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[30]), 
         .Z(delay_counter_31__N_531[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_853.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_854 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[29]), 
         .Z(delay_counter_31__N_531[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_854.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_855 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[28]), 
         .Z(delay_counter_31__N_531[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_855.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_856 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[27]), 
         .Z(delay_counter_31__N_531[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_856.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_857 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[26]), 
         .Z(delay_counter_31__N_531[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_857.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_858 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[25]), 
         .Z(delay_counter_31__N_531[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_858.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_859 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[24]), 
         .Z(delay_counter_31__N_531[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_859.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_860 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[23]), 
         .Z(delay_counter_31__N_531[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_860.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_861 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[22]), 
         .Z(delay_counter_31__N_531[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_861.init = 16'h2020;
    LUT4 i3_4_lut (.A(spi_byte_counter[0]), .B(spi_byte_counter[1]), .C(spi_byte_counter[2]), 
         .D(n131), .Z(n49273)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i3_4_lut.init = 16'h0800;
    LUT4 mux_129_i17_3_lut (.A(n2[23]), .B(DATA_OUT[0]), .C(n14326), .Z(WrData_23__N_691[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_862 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[21]), 
         .Z(delay_counter_31__N_531[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_862.init = 16'h2020;
    LUT4 mux_129_i18_3_lut (.A(n2[23]), .B(DATA_OUT[1]), .C(n14326), .Z(WrData_23__N_691[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i18_3_lut.init = 16'hcaca;
    LUT4 mux_129_i19_3_lut (.A(n2[23]), .B(DATA_OUT[2]), .C(n14326), .Z(WrData_23__N_691[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i19_3_lut.init = 16'hcaca;
    LUT4 mux_129_i20_3_lut (.A(n2[23]), .B(DATA_OUT[3]), .C(n14326), .Z(WrData_23__N_691[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i20_3_lut.init = 16'hcaca;
    LUT4 mux_129_i21_3_lut (.A(n2[23]), .B(DATA_OUT[4]), .C(n14326), .Z(WrData_23__N_691[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i21_3_lut.init = 16'hcaca;
    LUT4 mux_129_i22_3_lut (.A(n2[23]), .B(DATA_OUT[5]), .C(n14326), .Z(WrData_23__N_691[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i22_3_lut.init = 16'hcaca;
    LUT4 mux_129_i23_3_lut (.A(n2[23]), .B(DATA_OUT[6]), .C(n14326), .Z(WrData_23__N_691[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i23_3_lut.init = 16'hcaca;
    LUT4 mux_129_i24_3_lut (.A(n2[23]), .B(DATA_OUT[7]), .C(n14326), .Z(WrData_23__N_691[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i24_3_lut.init = 16'hcaca;
    LUT4 mux_143_i2_3_lut (.A(index[1]), .B(DATA_OUT[1]), .C(n14326), 
         .Z(WrAddr_8__N_747[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_863 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[20]), 
         .Z(delay_counter_31__N_531[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_863.init = 16'h2020;
    LUT4 mux_143_i3_3_lut (.A(index[2]), .B(DATA_OUT[2]), .C(n14326), 
         .Z(WrAddr_8__N_747[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i3_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_864 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[19]), 
         .Z(delay_counter_31__N_531[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_864.init = 16'h2020;
    LUT4 mux_143_i4_3_lut (.A(index[3]), .B(DATA_OUT[3]), .C(n14326), 
         .Z(WrAddr_8__N_747[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_865 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[18]), 
         .Z(delay_counter_31__N_531[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_865.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_866 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[17]), 
         .Z(delay_counter_31__N_531[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_866.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_867 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[16]), 
         .Z(delay_counter_31__N_531[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_867.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_868 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[15]), 
         .Z(delay_counter_31__N_531[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_868.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_869 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[14]), 
         .Z(delay_counter_31__N_531[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_869.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_870 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[13]), 
         .Z(delay_counter_31__N_531[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_870.init = 16'h2020;
    LUT4 mux_143_i5_3_lut (.A(index[4]), .B(DATA_OUT[4]), .C(n14326), 
         .Z(WrAddr_8__N_747[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_871 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[12]), 
         .Z(delay_counter_31__N_531[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_871.init = 16'h2020;
    LUT4 mux_143_i6_3_lut (.A(index[5]), .B(DATA_OUT[5]), .C(n14326), 
         .Z(WrAddr_8__N_747[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i6_3_lut.init = 16'hcaca;
    LUT4 mux_143_i7_3_lut (.A(index[6]), .B(DATA_OUT[6]), .C(n14326), 
         .Z(WrAddr_8__N_747[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i7_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_872 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[11]), 
         .Z(delay_counter_31__N_531[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_872.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_873 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[10]), 
         .Z(delay_counter_31__N_531[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_873.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_874 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[9]), 
         .Z(delay_counter_31__N_531[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_874.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_875 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[8]), 
         .Z(delay_counter_31__N_531[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_875.init = 16'h2020;
    PFUMX mux_206_Mux_2_i31 (.BLUT(n15), .ALUT(n50606), .C0(index[4]), 
          .Z(n2[23])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;
    LUT4 i1_2_lut_3_lut_adj_876 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[7]), 
         .Z(delay_counter_31__N_531[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_876.init = 16'h2020;
    LUT4 mux_143_i8_3_lut (.A(index[7]), .B(DATA_OUT[7]), .C(n14326), 
         .Z(WrAddr_8__N_747[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_877 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[6]), 
         .Z(delay_counter_31__N_531[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_877.init = 16'h2020;
    LUT4 mux_143_i9_3_lut (.A(index[8]), .B(DATA_OUT[0]), .C(n14326), 
         .Z(WrAddr_8__N_747[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_143_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_878 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[5]), 
         .Z(delay_counter_31__N_531[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_878.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_879 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[4]), 
         .Z(delay_counter_31__N_531[4])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_879.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_880 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[3]), 
         .Z(delay_counter_31__N_531[3])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_880.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_881 (.A(n55544), .B(n55545), .C(delay_counter_31__N_659[1]), 
         .Z(delay_counter_31__N_531[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i1_2_lut_3_lut_adj_881.init = 16'h2020;
    PFUMX i38895 (.BLUT(n54880), .ALUT(n54881), .C0(n14501), .Z(n54553));
    PFUMX mux_206_Mux_1_i31 (.BLUT(n15_adj_916), .ALUT(n30), .C0(index[4]), 
          .Z(n2[15])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;
    PFUMX mux_206_Mux_0_i31 (.BLUT(n15_adj_917), .ALUT(n50674), .C0(index[4]), 
          .Z(n2[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;
    CCU2D add_202_33 (.A0(index[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48210), 
          .S0(index_31__N_848[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_33.INIT0 = 16'h5aaa;
    defparam add_202_33.INIT1 = 16'h0000;
    defparam add_202_33.INJECT1_0 = "NO";
    defparam add_202_33.INJECT1_1 = "NO";
    CCU2D add_202_31 (.A0(index[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48209), .COUT(n48210), .S0(index_31__N_848[29]), .S1(index_31__N_848[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_31.INIT0 = 16'h5aaa;
    defparam add_202_31.INIT1 = 16'h5aaa;
    defparam add_202_31.INJECT1_0 = "NO";
    defparam add_202_31.INJECT1_1 = "NO";
    CCU2D add_202_29 (.A0(index[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48208), .COUT(n48209), .S0(index_31__N_848[27]), .S1(index_31__N_848[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_29.INIT0 = 16'h5aaa;
    defparam add_202_29.INIT1 = 16'h5aaa;
    defparam add_202_29.INJECT1_0 = "NO";
    defparam add_202_29.INJECT1_1 = "NO";
    CCU2D add_202_27 (.A0(index[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48207), .COUT(n48208), .S0(index_31__N_848[25]), .S1(index_31__N_848[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_27.INIT0 = 16'h5aaa;
    defparam add_202_27.INIT1 = 16'h5aaa;
    defparam add_202_27.INJECT1_0 = "NO";
    defparam add_202_27.INJECT1_1 = "NO";
    CCU2D add_202_25 (.A0(index[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48206), .COUT(n48207), .S0(index_31__N_848[23]), .S1(index_31__N_848[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_25.INIT0 = 16'h5aaa;
    defparam add_202_25.INIT1 = 16'h5aaa;
    defparam add_202_25.INJECT1_0 = "NO";
    defparam add_202_25.INJECT1_1 = "NO";
    CCU2D add_202_23 (.A0(index[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48205), .COUT(n48206), .S0(index_31__N_848[21]), .S1(index_31__N_848[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_23.INIT0 = 16'h5aaa;
    defparam add_202_23.INIT1 = 16'h5aaa;
    defparam add_202_23.INJECT1_0 = "NO";
    defparam add_202_23.INJECT1_1 = "NO";
    CCU2D add_202_21 (.A0(index[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48204), .COUT(n48205), .S0(index_31__N_848[19]), .S1(index_31__N_848[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_21.INIT0 = 16'h5aaa;
    defparam add_202_21.INIT1 = 16'h5aaa;
    defparam add_202_21.INJECT1_0 = "NO";
    defparam add_202_21.INJECT1_1 = "NO";
    CCU2D add_202_19 (.A0(index[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48203), .COUT(n48204), .S0(index_31__N_848[17]), .S1(index_31__N_848[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_19.INIT0 = 16'h5aaa;
    defparam add_202_19.INIT1 = 16'h5aaa;
    defparam add_202_19.INJECT1_0 = "NO";
    defparam add_202_19.INJECT1_1 = "NO";
    CCU2D add_202_17 (.A0(index[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48202), .COUT(n48203), .S0(index_31__N_848[15]), .S1(index_31__N_848[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_17.INIT0 = 16'h5aaa;
    defparam add_202_17.INIT1 = 16'h5aaa;
    defparam add_202_17.INJECT1_0 = "NO";
    defparam add_202_17.INJECT1_1 = "NO";
    CCU2D add_202_15 (.A0(index[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48201), .COUT(n48202), .S0(index_31__N_848[13]), .S1(index_31__N_848[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_15.INIT0 = 16'h5aaa;
    defparam add_202_15.INIT1 = 16'h5aaa;
    defparam add_202_15.INJECT1_0 = "NO";
    defparam add_202_15.INJECT1_1 = "NO";
    CCU2D add_202_13 (.A0(index[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48200), .COUT(n48201), .S0(index_31__N_848[11]), .S1(index_31__N_848[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_13.INIT0 = 16'h5aaa;
    defparam add_202_13.INIT1 = 16'h5aaa;
    defparam add_202_13.INJECT1_0 = "NO";
    defparam add_202_13.INJECT1_1 = "NO";
    CCU2D add_202_11 (.A0(index[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48199), .COUT(n48200), .S0(index_31__N_848[9]), .S1(index_31__N_848[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_11.INIT0 = 16'h5aaa;
    defparam add_202_11.INIT1 = 16'h5aaa;
    defparam add_202_11.INJECT1_0 = "NO";
    defparam add_202_11.INJECT1_1 = "NO";
    CCU2D add_202_9 (.A0(index[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48198), 
          .COUT(n48199), .S0(index_31__N_848[7]), .S1(index_31__N_848[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_9.INIT0 = 16'h5aaa;
    defparam add_202_9.INIT1 = 16'h5aaa;
    defparam add_202_9.INJECT1_0 = "NO";
    defparam add_202_9.INJECT1_1 = "NO";
    CCU2D add_202_7 (.A0(index[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48197), 
          .COUT(n48198), .S0(index_31__N_848[5]), .S1(index_31__N_848[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_7.INIT0 = 16'h5aaa;
    defparam add_202_7.INIT1 = 16'h5aaa;
    defparam add_202_7.INJECT1_0 = "NO";
    defparam add_202_7.INJECT1_1 = "NO";
    CCU2D add_202_5 (.A0(index[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48196), 
          .COUT(n48197), .S0(index_31__N_848[3]), .S1(index_31__N_848[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_5.INIT0 = 16'h5aaa;
    defparam add_202_5.INIT1 = 16'h5aaa;
    defparam add_202_5.INJECT1_0 = "NO";
    defparam add_202_5.INJECT1_1 = "NO";
    CCU2D add_33925_32 (.A0(spi_byte_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n49038), .S1(n14361));
    defparam add_33925_32.INIT0 = 16'hf555;
    defparam add_33925_32.INIT1 = 16'h0000;
    defparam add_33925_32.INJECT1_0 = "NO";
    defparam add_33925_32.INJECT1_1 = "NO";
    CCU2D add_33925_30 (.A0(spi_byte_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49037), .COUT(n49038));
    defparam add_33925_30.INIT0 = 16'h5555;
    defparam add_33925_30.INIT1 = 16'h5555;
    defparam add_33925_30.INJECT1_0 = "NO";
    defparam add_33925_30.INJECT1_1 = "NO";
    LUT4 mux_132_i5_3_lut (.A(index[4]), .B(DATA_OUT[5]), .C(n14326), 
         .Z(fb_31__N_715[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_132_i5_3_lut.init = 16'hcaca;
    CCU2D add_33925_28 (.A0(spi_byte_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49036), .COUT(n49037));
    defparam add_33925_28.INIT0 = 16'h5555;
    defparam add_33925_28.INIT1 = 16'h5555;
    defparam add_33925_28.INJECT1_0 = "NO";
    defparam add_33925_28.INJECT1_1 = "NO";
    CCU2D add_33925_26 (.A0(spi_byte_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49035), .COUT(n49036));
    defparam add_33925_26.INIT0 = 16'h5555;
    defparam add_33925_26.INIT1 = 16'h5555;
    defparam add_33925_26.INJECT1_0 = "NO";
    defparam add_33925_26.INJECT1_1 = "NO";
    CCU2D add_33925_24 (.A0(spi_byte_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49034), .COUT(n49035));
    defparam add_33925_24.INIT0 = 16'h5555;
    defparam add_33925_24.INIT1 = 16'h5555;
    defparam add_33925_24.INJECT1_0 = "NO";
    defparam add_33925_24.INJECT1_1 = "NO";
    CCU2D add_33925_22 (.A0(spi_byte_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49033), .COUT(n49034));
    defparam add_33925_22.INIT0 = 16'h5555;
    defparam add_33925_22.INIT1 = 16'h5555;
    defparam add_33925_22.INJECT1_0 = "NO";
    defparam add_33925_22.INJECT1_1 = "NO";
    CCU2D add_33925_20 (.A0(spi_byte_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49032), .COUT(n49033));
    defparam add_33925_20.INIT0 = 16'h5555;
    defparam add_33925_20.INIT1 = 16'h5555;
    defparam add_33925_20.INJECT1_0 = "NO";
    defparam add_33925_20.INJECT1_1 = "NO";
    CCU2D add_33925_18 (.A0(spi_byte_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49031), .COUT(n49032));
    defparam add_33925_18.INIT0 = 16'h5555;
    defparam add_33925_18.INIT1 = 16'h5555;
    defparam add_33925_18.INJECT1_0 = "NO";
    defparam add_33925_18.INJECT1_1 = "NO";
    CCU2D add_202_3 (.A0(index[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48195), 
          .COUT(n48196), .S0(index_31__N_848[1]), .S1(index_31__N_848[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_3.INIT0 = 16'h5aaa;
    defparam add_202_3.INIT1 = 16'h5aaa;
    defparam add_202_3.INJECT1_0 = "NO";
    defparam add_202_3.INJECT1_1 = "NO";
    CCU2D add_33925_16 (.A0(spi_byte_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49030), .COUT(n49031));
    defparam add_33925_16.INIT0 = 16'h5555;
    defparam add_33925_16.INIT1 = 16'h5555;
    defparam add_33925_16.INJECT1_0 = "NO";
    defparam add_33925_16.INJECT1_1 = "NO";
    CCU2D add_33925_14 (.A0(spi_byte_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49029), .COUT(n49030));
    defparam add_33925_14.INIT0 = 16'h5555;
    defparam add_33925_14.INIT1 = 16'h5555;
    defparam add_33925_14.INJECT1_0 = "NO";
    defparam add_33925_14.INJECT1_1 = "NO";
    CCU2D add_202_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[0]), .B1(n14326), .C1(GND_net), .D1(GND_net), .COUT(n48195), 
          .S1(index_31__N_848[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(110[15:20])
    defparam add_202_1.INIT0 = 16'hF000;
    defparam add_202_1.INIT1 = 16'h5999;
    defparam add_202_1.INJECT1_0 = "NO";
    defparam add_202_1.INJECT1_1 = "NO";
    CCU2D add_33925_12 (.A0(spi_byte_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49028), .COUT(n49029));
    defparam add_33925_12.INIT0 = 16'h5555;
    defparam add_33925_12.INIT1 = 16'h5555;
    defparam add_33925_12.INJECT1_0 = "NO";
    defparam add_33925_12.INJECT1_1 = "NO";
    CCU2D add_33925_10 (.A0(spi_byte_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49027), .COUT(n49028));
    defparam add_33925_10.INIT0 = 16'h5555;
    defparam add_33925_10.INIT1 = 16'h5555;
    defparam add_33925_10.INJECT1_0 = "NO";
    defparam add_33925_10.INJECT1_1 = "NO";
    CCU2D add_33925_8 (.A0(spi_byte_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49026), .COUT(n49027));
    defparam add_33925_8.INIT0 = 16'h5555;
    defparam add_33925_8.INIT1 = 16'h5555;
    defparam add_33925_8.INJECT1_0 = "NO";
    defparam add_33925_8.INJECT1_1 = "NO";
    CCU2D add_33925_6 (.A0(spi_byte_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49025), .COUT(n49026));
    defparam add_33925_6.INIT0 = 16'h5555;
    defparam add_33925_6.INIT1 = 16'h5555;
    defparam add_33925_6.INJECT1_0 = "NO";
    defparam add_33925_6.INJECT1_1 = "NO";
    CCU2D add_33925_4 (.A0(spi_byte_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49024), .COUT(n49025));
    defparam add_33925_4.INIT0 = 16'h5555;
    defparam add_33925_4.INIT1 = 16'h5555;
    defparam add_33925_4.INJECT1_0 = "NO";
    defparam add_33925_4.INJECT1_1 = "NO";
    CCU2D add_33925_2 (.A0(spi_byte_counter[1]), .B0(spi_byte_counter[0]), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n49024));
    defparam add_33925_2.INIT0 = 16'h1000;
    defparam add_33925_2.INIT1 = 16'h5555;
    defparam add_33925_2.INJECT1_0 = "NO";
    defparam add_33925_2.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(n14396), .B(n14326), .C(n54679), .D(n54741), 
         .Z(sclk_c_enable_1284)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h7300;
    CCU2D add_123_33 (.A0(spi_byte_timeout[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48194), .S0(n869[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_33.INIT0 = 16'h5555;
    defparam add_123_33.INIT1 = 16'h0000;
    defparam add_123_33.INJECT1_0 = "NO";
    defparam add_123_33.INJECT1_1 = "NO";
    CCU2D add_123_31 (.A0(spi_byte_timeout[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48193), .COUT(n48194), .S0(n869[29]), 
          .S1(n869[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_31.INIT0 = 16'h5555;
    defparam add_123_31.INIT1 = 16'h5555;
    defparam add_123_31.INJECT1_0 = "NO";
    defparam add_123_31.INJECT1_1 = "NO";
    CCU2D add_123_29 (.A0(spi_byte_timeout[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48192), .COUT(n48193), .S0(n869[27]), 
          .S1(n869[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_29.INIT0 = 16'h5555;
    defparam add_123_29.INIT1 = 16'h5555;
    defparam add_123_29.INJECT1_0 = "NO";
    defparam add_123_29.INJECT1_1 = "NO";
    CCU2D add_123_27 (.A0(spi_byte_timeout[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48191), .COUT(n48192), .S0(n869[25]), 
          .S1(n869[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_27.INIT0 = 16'h5555;
    defparam add_123_27.INIT1 = 16'h5555;
    defparam add_123_27.INJECT1_0 = "NO";
    defparam add_123_27.INJECT1_1 = "NO";
    CCU2D add_123_25 (.A0(spi_byte_timeout[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48190), .COUT(n48191), .S0(n869[23]), 
          .S1(n869[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_25.INIT0 = 16'h5555;
    defparam add_123_25.INIT1 = 16'h5555;
    defparam add_123_25.INJECT1_0 = "NO";
    defparam add_123_25.INJECT1_1 = "NO";
    CCU2D add_123_23 (.A0(spi_byte_timeout[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48189), .COUT(n48190), .S0(n869[21]), 
          .S1(n869[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_23.INIT0 = 16'h5555;
    defparam add_123_23.INIT1 = 16'h5555;
    defparam add_123_23.INJECT1_0 = "NO";
    defparam add_123_23.INJECT1_1 = "NO";
    CCU2D add_123_21 (.A0(spi_byte_timeout[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48188), .COUT(n48189), .S0(n869[19]), 
          .S1(n869[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_21.INIT0 = 16'h5555;
    defparam add_123_21.INIT1 = 16'h5555;
    defparam add_123_21.INJECT1_0 = "NO";
    defparam add_123_21.INJECT1_1 = "NO";
    CCU2D add_123_19 (.A0(spi_byte_timeout[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48187), .COUT(n48188), .S0(n869[17]), 
          .S1(n869[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_19.INIT0 = 16'h5555;
    defparam add_123_19.INIT1 = 16'h5555;
    defparam add_123_19.INJECT1_0 = "NO";
    defparam add_123_19.INJECT1_1 = "NO";
    CCU2D add_123_17 (.A0(spi_byte_timeout[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48186), .COUT(n48187), .S0(n869[15]), 
          .S1(n869[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_17.INIT0 = 16'h5555;
    defparam add_123_17.INIT1 = 16'h5555;
    defparam add_123_17.INJECT1_0 = "NO";
    defparam add_123_17.INJECT1_1 = "NO";
    CCU2D add_123_15 (.A0(spi_byte_timeout[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48185), .COUT(n48186), .S0(n869[13]), 
          .S1(n869[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_15.INIT0 = 16'h5555;
    defparam add_123_15.INIT1 = 16'h5555;
    defparam add_123_15.INJECT1_0 = "NO";
    defparam add_123_15.INJECT1_1 = "NO";
    CCU2D add_123_13 (.A0(spi_byte_timeout[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48184), .COUT(n48185), .S0(n869[11]), 
          .S1(n869[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_13.INIT0 = 16'h5555;
    defparam add_123_13.INIT1 = 16'h5555;
    defparam add_123_13.INJECT1_0 = "NO";
    defparam add_123_13.INJECT1_1 = "NO";
    CCU2D add_123_11 (.A0(spi_byte_timeout[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48183), .COUT(n48184), .S0(n869[9]), .S1(n869[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_11.INIT0 = 16'h5555;
    defparam add_123_11.INIT1 = 16'h5555;
    defparam add_123_11.INJECT1_0 = "NO";
    defparam add_123_11.INJECT1_1 = "NO";
    CCU2D add_123_9 (.A0(spi_byte_timeout[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48182), .COUT(n48183), .S0(n869[7]), .S1(n869[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_9.INIT0 = 16'h5555;
    defparam add_123_9.INIT1 = 16'h5555;
    defparam add_123_9.INJECT1_0 = "NO";
    defparam add_123_9.INJECT1_1 = "NO";
    CCU2D add_123_7 (.A0(spi_byte_timeout[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48181), .COUT(n48182), .S0(n869[5]), .S1(n869[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_7.INIT0 = 16'h5555;
    defparam add_123_7.INIT1 = 16'h5555;
    defparam add_123_7.INJECT1_0 = "NO";
    defparam add_123_7.INJECT1_1 = "NO";
    CCU2D add_33927_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48991), 
          .S0(n14571));
    defparam add_33927_cout.INIT0 = 16'h0000;
    defparam add_33927_cout.INIT1 = 16'h0000;
    defparam add_33927_cout.INJECT1_0 = "NO";
    defparam add_33927_cout.INJECT1_1 = "NO";
    CCU2D add_33927_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48990), .COUT(n48991));
    defparam add_33927_31.INIT0 = 16'hf555;
    defparam add_33927_31.INIT1 = 16'h5555;
    defparam add_33927_31.INJECT1_0 = "NO";
    defparam add_33927_31.INJECT1_1 = "NO";
    CCU2D add_33927_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48989), .COUT(n48990));
    defparam add_33927_29.INIT0 = 16'hf555;
    defparam add_33927_29.INIT1 = 16'hf555;
    defparam add_33927_29.INJECT1_0 = "NO";
    defparam add_33927_29.INJECT1_1 = "NO";
    CCU2D add_33927_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48988), .COUT(n48989));
    defparam add_33927_27.INIT0 = 16'hf555;
    defparam add_33927_27.INIT1 = 16'hf555;
    defparam add_33927_27.INJECT1_0 = "NO";
    defparam add_33927_27.INJECT1_1 = "NO";
    CCU2D add_33927_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48987), .COUT(n48988));
    defparam add_33927_25.INIT0 = 16'hf555;
    defparam add_33927_25.INIT1 = 16'hf555;
    defparam add_33927_25.INJECT1_0 = "NO";
    defparam add_33927_25.INJECT1_1 = "NO";
    CCU2D add_33927_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48986), .COUT(n48987));
    defparam add_33927_23.INIT0 = 16'hf555;
    defparam add_33927_23.INIT1 = 16'hf555;
    defparam add_33927_23.INJECT1_0 = "NO";
    defparam add_33927_23.INJECT1_1 = "NO";
    CCU2D add_33927_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48985), .COUT(n48986));
    defparam add_33927_21.INIT0 = 16'hf555;
    defparam add_33927_21.INIT1 = 16'hf555;
    defparam add_33927_21.INJECT1_0 = "NO";
    defparam add_33927_21.INJECT1_1 = "NO";
    CCU2D add_33927_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48984), .COUT(n48985));
    defparam add_33927_19.INIT0 = 16'hf555;
    defparam add_33927_19.INIT1 = 16'hf555;
    defparam add_33927_19.INJECT1_0 = "NO";
    defparam add_33927_19.INJECT1_1 = "NO";
    CCU2D add_33927_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48983), .COUT(n48984));
    defparam add_33927_17.INIT0 = 16'hf555;
    defparam add_33927_17.INIT1 = 16'hf555;
    defparam add_33927_17.INJECT1_0 = "NO";
    defparam add_33927_17.INJECT1_1 = "NO";
    CCU2D add_33927_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48982), .COUT(n48983));
    defparam add_33927_15.INIT0 = 16'hf555;
    defparam add_33927_15.INIT1 = 16'hf555;
    defparam add_33927_15.INJECT1_0 = "NO";
    defparam add_33927_15.INJECT1_1 = "NO";
    CCU2D add_33927_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48981), .COUT(n48982));
    defparam add_33927_13.INIT0 = 16'hf555;
    defparam add_33927_13.INIT1 = 16'hf555;
    defparam add_33927_13.INJECT1_0 = "NO";
    defparam add_33927_13.INJECT1_1 = "NO";
    CCU2D add_33927_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48980), .COUT(n48981));
    defparam add_33927_11.INIT0 = 16'hf555;
    defparam add_33927_11.INIT1 = 16'hf555;
    defparam add_33927_11.INJECT1_0 = "NO";
    defparam add_33927_11.INJECT1_1 = "NO";
    CCU2D add_33927_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48979), .COUT(n48980));
    defparam add_33927_9.INIT0 = 16'hf555;
    defparam add_33927_9.INIT1 = 16'hf555;
    defparam add_33927_9.INJECT1_0 = "NO";
    defparam add_33927_9.INJECT1_1 = "NO";
    CCU2D add_123_5 (.A0(spi_byte_timeout[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48180), .COUT(n48181), .S0(n869[3]), .S1(n869[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_5.INIT0 = 16'h5555;
    defparam add_123_5.INIT1 = 16'h5555;
    defparam add_123_5.INJECT1_0 = "NO";
    defparam add_123_5.INJECT1_1 = "NO";
    CCU2D add_33927_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48978), .COUT(n48979));
    defparam add_33927_7.INIT0 = 16'hf555;
    defparam add_33927_7.INIT1 = 16'hf555;
    defparam add_33927_7.INJECT1_0 = "NO";
    defparam add_33927_7.INJECT1_1 = "NO";
    CCU2D add_33927_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48977), .COUT(n48978));
    defparam add_33927_5.INIT0 = 16'hf555;
    defparam add_33927_5.INIT1 = 16'hf555;
    defparam add_33927_5.INJECT1_0 = "NO";
    defparam add_33927_5.INJECT1_1 = "NO";
    CCU2D add_33927_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48976), .COUT(n48977));
    defparam add_33927_3.INIT0 = 16'hf555;
    defparam add_33927_3.INIT1 = 16'hf555;
    defparam add_33927_3.INJECT1_0 = "NO";
    defparam add_33927_3.INJECT1_1 = "NO";
    CCU2D add_33927_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48976));
    defparam add_33927_1.INIT0 = 16'hF000;
    defparam add_33927_1.INIT1 = 16'ha666;
    defparam add_33927_1.INJECT1_0 = "NO";
    defparam add_33927_1.INJECT1_1 = "NO";
    CCU2D add_33928_30 (.A0(index[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48975), 
          .S1(n14326));
    defparam add_33928_30.INIT0 = 16'hf555;
    defparam add_33928_30.INIT1 = 16'h0000;
    defparam add_33928_30.INJECT1_0 = "NO";
    defparam add_33928_30.INJECT1_1 = "NO";
    CCU2D add_33928_28 (.A0(index[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48974), .COUT(n48975));
    defparam add_33928_28.INIT0 = 16'h5555;
    defparam add_33928_28.INIT1 = 16'h5555;
    defparam add_33928_28.INJECT1_0 = "NO";
    defparam add_33928_28.INJECT1_1 = "NO";
    CCU2D add_33928_26 (.A0(index[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48973), .COUT(n48974));
    defparam add_33928_26.INIT0 = 16'h5555;
    defparam add_33928_26.INIT1 = 16'h5555;
    defparam add_33928_26.INJECT1_0 = "NO";
    defparam add_33928_26.INJECT1_1 = "NO";
    CCU2D add_33928_24 (.A0(index[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48972), .COUT(n48973));
    defparam add_33928_24.INIT0 = 16'h5555;
    defparam add_33928_24.INIT1 = 16'h5555;
    defparam add_33928_24.INJECT1_0 = "NO";
    defparam add_33928_24.INJECT1_1 = "NO";
    CCU2D add_33928_22 (.A0(index[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48971), .COUT(n48972));
    defparam add_33928_22.INIT0 = 16'h5555;
    defparam add_33928_22.INIT1 = 16'h5555;
    defparam add_33928_22.INJECT1_0 = "NO";
    defparam add_33928_22.INJECT1_1 = "NO";
    CCU2D add_33928_20 (.A0(index[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48970), .COUT(n48971));
    defparam add_33928_20.INIT0 = 16'h5555;
    defparam add_33928_20.INIT1 = 16'h5555;
    defparam add_33928_20.INJECT1_0 = "NO";
    defparam add_33928_20.INJECT1_1 = "NO";
    CCU2D add_33928_18 (.A0(index[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48969), .COUT(n48970));
    defparam add_33928_18.INIT0 = 16'h5555;
    defparam add_33928_18.INIT1 = 16'h5555;
    defparam add_33928_18.INJECT1_0 = "NO";
    defparam add_33928_18.INJECT1_1 = "NO";
    CCU2D add_33928_16 (.A0(index[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48968), .COUT(n48969));
    defparam add_33928_16.INIT0 = 16'h5555;
    defparam add_33928_16.INIT1 = 16'h5555;
    defparam add_33928_16.INJECT1_0 = "NO";
    defparam add_33928_16.INJECT1_1 = "NO";
    CCU2D add_33928_14 (.A0(index[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48967), .COUT(n48968));
    defparam add_33928_14.INIT0 = 16'h5555;
    defparam add_33928_14.INIT1 = 16'h5555;
    defparam add_33928_14.INJECT1_0 = "NO";
    defparam add_33928_14.INJECT1_1 = "NO";
    CCU2D add_123_3 (.A0(spi_byte_timeout[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_timeout[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48179), .COUT(n48180), .S0(n869[1]), .S1(n869[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_3.INIT0 = 16'h5555;
    defparam add_123_3.INIT1 = 16'h5555;
    defparam add_123_3.INJECT1_0 = "NO";
    defparam add_123_3.INJECT1_1 = "NO";
    CCU2D add_123_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(spi_byte_timeout[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48179), .S1(n869[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(82[26:42])
    defparam add_123_1.INIT0 = 16'hF000;
    defparam add_123_1.INIT1 = 16'h5555;
    defparam add_123_1.INJECT1_0 = "NO";
    defparam add_123_1.INJECT1_1 = "NO";
    CCU2D add_117_33 (.A0(spi_byte_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48178), .S0(n830[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_33.INIT0 = 16'h5aaa;
    defparam add_117_33.INIT1 = 16'h0000;
    defparam add_117_33.INJECT1_0 = "NO";
    defparam add_117_33.INJECT1_1 = "NO";
    CCU2D add_117_31 (.A0(spi_byte_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48177), .COUT(n48178), .S0(n830[29]), 
          .S1(n830[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_31.INIT0 = 16'h5aaa;
    defparam add_117_31.INIT1 = 16'h5aaa;
    defparam add_117_31.INJECT1_0 = "NO";
    defparam add_117_31.INJECT1_1 = "NO";
    CCU2D add_117_29 (.A0(spi_byte_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48176), .COUT(n48177), .S0(n830[27]), 
          .S1(n830[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_29.INIT0 = 16'h5aaa;
    defparam add_117_29.INIT1 = 16'h5aaa;
    defparam add_117_29.INJECT1_0 = "NO";
    defparam add_117_29.INJECT1_1 = "NO";
    CCU2D add_117_27 (.A0(spi_byte_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48175), .COUT(n48176), .S0(n830[25]), 
          .S1(n830[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_27.INIT0 = 16'h5aaa;
    defparam add_117_27.INIT1 = 16'h5aaa;
    defparam add_117_27.INJECT1_0 = "NO";
    defparam add_117_27.INJECT1_1 = "NO";
    CCU2D add_117_25 (.A0(spi_byte_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48174), .COUT(n48175), .S0(n830[23]), 
          .S1(n830[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_25.INIT0 = 16'h5aaa;
    defparam add_117_25.INIT1 = 16'h5aaa;
    defparam add_117_25.INJECT1_0 = "NO";
    defparam add_117_25.INJECT1_1 = "NO";
    CCU2D add_117_23 (.A0(spi_byte_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48173), .COUT(n48174), .S0(n830[21]), 
          .S1(n830[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_23.INIT0 = 16'h5aaa;
    defparam add_117_23.INIT1 = 16'h5aaa;
    defparam add_117_23.INJECT1_0 = "NO";
    defparam add_117_23.INJECT1_1 = "NO";
    CCU2D add_33928_12 (.A0(index[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48966), .COUT(n48967));
    defparam add_33928_12.INIT0 = 16'h5555;
    defparam add_33928_12.INIT1 = 16'h5555;
    defparam add_33928_12.INJECT1_0 = "NO";
    defparam add_33928_12.INJECT1_1 = "NO";
    CCU2D add_117_21 (.A0(spi_byte_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48172), .COUT(n48173), .S0(n830[19]), 
          .S1(n830[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_21.INIT0 = 16'h5aaa;
    defparam add_117_21.INIT1 = 16'h5aaa;
    defparam add_117_21.INJECT1_0 = "NO";
    defparam add_117_21.INJECT1_1 = "NO";
    CCU2D add_117_19 (.A0(spi_byte_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48171), .COUT(n48172), .S0(n830[17]), 
          .S1(n830[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_19.INIT0 = 16'h5aaa;
    defparam add_117_19.INIT1 = 16'h5aaa;
    defparam add_117_19.INJECT1_0 = "NO";
    defparam add_117_19.INJECT1_1 = "NO";
    CCU2D add_117_17 (.A0(spi_byte_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48170), .COUT(n48171), .S0(n830[15]), 
          .S1(n830[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_17.INIT0 = 16'h5aaa;
    defparam add_117_17.INIT1 = 16'h5aaa;
    defparam add_117_17.INJECT1_0 = "NO";
    defparam add_117_17.INJECT1_1 = "NO";
    CCU2D add_117_15 (.A0(spi_byte_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48169), .COUT(n48170), .S0(n830[13]), 
          .S1(n830[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_15.INIT0 = 16'h5aaa;
    defparam add_117_15.INIT1 = 16'h5aaa;
    defparam add_117_15.INJECT1_0 = "NO";
    defparam add_117_15.INJECT1_1 = "NO";
    CCU2D add_117_13 (.A0(spi_byte_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48168), .COUT(n48169), .S0(n830[11]), 
          .S1(n830[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_13.INIT0 = 16'h5aaa;
    defparam add_117_13.INIT1 = 16'h5aaa;
    defparam add_117_13.INJECT1_0 = "NO";
    defparam add_117_13.INJECT1_1 = "NO";
    CCU2D add_33928_10 (.A0(index[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48965), .COUT(n48966));
    defparam add_33928_10.INIT0 = 16'h5555;
    defparam add_33928_10.INIT1 = 16'h5555;
    defparam add_33928_10.INJECT1_0 = "NO";
    defparam add_33928_10.INJECT1_1 = "NO";
    CCU2D add_33928_8 (.A0(index[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48964), .COUT(n48965));
    defparam add_33928_8.INIT0 = 16'h5555;
    defparam add_33928_8.INIT1 = 16'h5555;
    defparam add_33928_8.INJECT1_0 = "NO";
    defparam add_33928_8.INJECT1_1 = "NO";
    CCU2D add_33928_6 (.A0(index[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48963), 
          .COUT(n48964));
    defparam add_33928_6.INIT0 = 16'h5555;
    defparam add_33928_6.INIT1 = 16'h5555;
    defparam add_33928_6.INJECT1_0 = "NO";
    defparam add_33928_6.INJECT1_1 = "NO";
    CCU2D add_117_11 (.A0(spi_byte_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48167), .COUT(n48168), .S0(n830[9]), .S1(n830[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_11.INIT0 = 16'h5aaa;
    defparam add_117_11.INIT1 = 16'h5aaa;
    defparam add_117_11.INJECT1_0 = "NO";
    defparam add_117_11.INJECT1_1 = "NO";
    CCU2D add_117_9 (.A0(spi_byte_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48166), .COUT(n48167), .S0(n830[7]), .S1(n830[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_9.INIT0 = 16'h5aaa;
    defparam add_117_9.INIT1 = 16'h5aaa;
    defparam add_117_9.INJECT1_0 = "NO";
    defparam add_117_9.INJECT1_1 = "NO";
    CCU2D add_117_7 (.A0(spi_byte_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48165), .COUT(n48166), .S0(n830[5]), .S1(n830[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_7.INIT0 = 16'h5aaa;
    defparam add_117_7.INIT1 = 16'h5aaa;
    defparam add_117_7.INJECT1_0 = "NO";
    defparam add_117_7.INJECT1_1 = "NO";
    CCU2D add_117_5 (.A0(spi_byte_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48164), .COUT(n48165), .S0(n830[3]), .S1(n830[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_5.INIT0 = 16'h5aaa;
    defparam add_117_5.INIT1 = 16'h5aaa;
    defparam add_117_5.INJECT1_0 = "NO";
    defparam add_117_5.INJECT1_1 = "NO";
    CCU2D add_33928_4 (.A0(index[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(index[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48962), 
          .COUT(n48963));
    defparam add_33928_4.INIT0 = 16'h5555;
    defparam add_33928_4.INIT1 = 16'h5555;
    defparam add_33928_4.INJECT1_0 = "NO";
    defparam add_33928_4.INJECT1_1 = "NO";
    CCU2D add_117_3 (.A0(spi_byte_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48163), .COUT(n48164), .S0(n830[1]), .S1(n830[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_3.INIT0 = 16'h5aaa;
    defparam add_117_3.INIT1 = 16'h5aaa;
    defparam add_117_3.INJECT1_0 = "NO";
    defparam add_117_3.INJECT1_1 = "NO";
    CCU2D add_117_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(spi_byte_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48163), .S1(n830[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(79[26:42])
    defparam add_117_1.INIT0 = 16'hF000;
    defparam add_117_1.INIT1 = 16'h5555;
    defparam add_117_1.INJECT1_0 = "NO";
    defparam add_117_1.INJECT1_1 = "NO";
    CCU2D add_33928_2 (.A0(index[3]), .B0(index[2]), .C0(GND_net), .D0(GND_net), 
          .A1(index[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n48962));
    defparam add_33928_2.INIT0 = 16'h1000;
    defparam add_33928_2.INIT1 = 16'h5aaa;
    defparam add_33928_2.INJECT1_0 = "NO";
    defparam add_33928_2.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47914), .S0(n14396));
    defparam sub_3233_add_2_cout.INIT0 = 16'h0000;
    defparam sub_3233_add_2_cout.INIT1 = 16'h0000;
    defparam sub_3233_add_2_cout.INJECT1_0 = "NO";
    defparam sub_3233_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_32 (.A0(spi_byte_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47913), .COUT(n47914));
    defparam sub_3233_add_2_32.INIT0 = 16'h5555;
    defparam sub_3233_add_2_32.INIT1 = 16'hf555;
    defparam sub_3233_add_2_32.INJECT1_0 = "NO";
    defparam sub_3233_add_2_32.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_30 (.A0(spi_byte_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47912), .COUT(n47913));
    defparam sub_3233_add_2_30.INIT0 = 16'h5555;
    defparam sub_3233_add_2_30.INIT1 = 16'h5555;
    defparam sub_3233_add_2_30.INJECT1_0 = "NO";
    defparam sub_3233_add_2_30.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_28 (.A0(spi_byte_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47911), .COUT(n47912));
    defparam sub_3233_add_2_28.INIT0 = 16'h5555;
    defparam sub_3233_add_2_28.INIT1 = 16'h5555;
    defparam sub_3233_add_2_28.INJECT1_0 = "NO";
    defparam sub_3233_add_2_28.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_26 (.A0(spi_byte_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47910), .COUT(n47911));
    defparam sub_3233_add_2_26.INIT0 = 16'h5555;
    defparam sub_3233_add_2_26.INIT1 = 16'h5555;
    defparam sub_3233_add_2_26.INJECT1_0 = "NO";
    defparam sub_3233_add_2_26.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_24 (.A0(spi_byte_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47909), .COUT(n47910));
    defparam sub_3233_add_2_24.INIT0 = 16'h5555;
    defparam sub_3233_add_2_24.INIT1 = 16'h5555;
    defparam sub_3233_add_2_24.INJECT1_0 = "NO";
    defparam sub_3233_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_22 (.A0(spi_byte_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47908), .COUT(n47909));
    defparam sub_3233_add_2_22.INIT0 = 16'h5555;
    defparam sub_3233_add_2_22.INIT1 = 16'h5555;
    defparam sub_3233_add_2_22.INJECT1_0 = "NO";
    defparam sub_3233_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_20 (.A0(spi_byte_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47907), .COUT(n47908));
    defparam sub_3233_add_2_20.INIT0 = 16'h5555;
    defparam sub_3233_add_2_20.INIT1 = 16'h5555;
    defparam sub_3233_add_2_20.INJECT1_0 = "NO";
    defparam sub_3233_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_18 (.A0(spi_byte_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47906), .COUT(n47907));
    defparam sub_3233_add_2_18.INIT0 = 16'h5555;
    defparam sub_3233_add_2_18.INIT1 = 16'h5555;
    defparam sub_3233_add_2_18.INJECT1_0 = "NO";
    defparam sub_3233_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_16 (.A0(spi_byte_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47905), .COUT(n47906));
    defparam sub_3233_add_2_16.INIT0 = 16'h5555;
    defparam sub_3233_add_2_16.INIT1 = 16'h5555;
    defparam sub_3233_add_2_16.INJECT1_0 = "NO";
    defparam sub_3233_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_14 (.A0(spi_byte_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47904), .COUT(n47905));
    defparam sub_3233_add_2_14.INIT0 = 16'h5555;
    defparam sub_3233_add_2_14.INIT1 = 16'h5555;
    defparam sub_3233_add_2_14.INJECT1_0 = "NO";
    defparam sub_3233_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_12 (.A0(spi_byte_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47903), .COUT(n47904));
    defparam sub_3233_add_2_12.INIT0 = 16'h5555;
    defparam sub_3233_add_2_12.INIT1 = 16'h5555;
    defparam sub_3233_add_2_12.INJECT1_0 = "NO";
    defparam sub_3233_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_10 (.A0(spi_byte_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47902), .COUT(n47903));
    defparam sub_3233_add_2_10.INIT0 = 16'h5555;
    defparam sub_3233_add_2_10.INIT1 = 16'h5555;
    defparam sub_3233_add_2_10.INJECT1_0 = "NO";
    defparam sub_3233_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_8 (.A0(spi_byte_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47901), .COUT(n47902));
    defparam sub_3233_add_2_8.INIT0 = 16'h5555;
    defparam sub_3233_add_2_8.INIT1 = 16'h5555;
    defparam sub_3233_add_2_8.INJECT1_0 = "NO";
    defparam sub_3233_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_6 (.A0(spi_byte_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47900), .COUT(n47901));
    defparam sub_3233_add_2_6.INIT0 = 16'h5555;
    defparam sub_3233_add_2_6.INIT1 = 16'h5555;
    defparam sub_3233_add_2_6.INJECT1_0 = "NO";
    defparam sub_3233_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_4 (.A0(spi_byte_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47899), .COUT(n47900));
    defparam sub_3233_add_2_4.INIT0 = 16'h5555;
    defparam sub_3233_add_2_4.INIT1 = 16'h5555;
    defparam sub_3233_add_2_4.INJECT1_0 = "NO";
    defparam sub_3233_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_3233_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[1]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n47899));
    defparam sub_3233_add_2_2.INIT0 = 16'h0000;
    defparam sub_3233_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_3233_add_2_2.INJECT1_0 = "NO";
    defparam sub_3233_add_2_2.INJECT1_1 = "NO";
    CCU2D add_33918_32 (.A0(spi_byte_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48417), .S1(n14431));
    defparam add_33918_32.INIT0 = 16'hf555;
    defparam add_33918_32.INIT1 = 16'h0000;
    defparam add_33918_32.INJECT1_0 = "NO";
    defparam add_33918_32.INJECT1_1 = "NO";
    CCU2D add_33918_30 (.A0(spi_byte_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48416), .COUT(n48417));
    defparam add_33918_30.INIT0 = 16'h5555;
    defparam add_33918_30.INIT1 = 16'h5555;
    defparam add_33918_30.INJECT1_0 = "NO";
    defparam add_33918_30.INJECT1_1 = "NO";
    CCU2D add_33918_28 (.A0(spi_byte_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48415), .COUT(n48416));
    defparam add_33918_28.INIT0 = 16'h5555;
    defparam add_33918_28.INIT1 = 16'h5555;
    defparam add_33918_28.INJECT1_0 = "NO";
    defparam add_33918_28.INJECT1_1 = "NO";
    CCU2D add_33918_26 (.A0(spi_byte_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48414), .COUT(n48415));
    defparam add_33918_26.INIT0 = 16'h5555;
    defparam add_33918_26.INIT1 = 16'h5555;
    defparam add_33918_26.INJECT1_0 = "NO";
    defparam add_33918_26.INJECT1_1 = "NO";
    CCU2D add_33918_24 (.A0(spi_byte_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48413), .COUT(n48414));
    defparam add_33918_24.INIT0 = 16'h5555;
    defparam add_33918_24.INIT1 = 16'h5555;
    defparam add_33918_24.INJECT1_0 = "NO";
    defparam add_33918_24.INJECT1_1 = "NO";
    CCU2D add_33918_22 (.A0(spi_byte_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48412), .COUT(n48413));
    defparam add_33918_22.INIT0 = 16'h5555;
    defparam add_33918_22.INIT1 = 16'h5555;
    defparam add_33918_22.INJECT1_0 = "NO";
    defparam add_33918_22.INJECT1_1 = "NO";
    CCU2D add_33918_20 (.A0(spi_byte_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48411), .COUT(n48412));
    defparam add_33918_20.INIT0 = 16'h5555;
    defparam add_33918_20.INIT1 = 16'h5555;
    defparam add_33918_20.INJECT1_0 = "NO";
    defparam add_33918_20.INJECT1_1 = "NO";
    CCU2D add_33918_18 (.A0(spi_byte_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48410), .COUT(n48411));
    defparam add_33918_18.INIT0 = 16'h5555;
    defparam add_33918_18.INIT1 = 16'h5555;
    defparam add_33918_18.INJECT1_0 = "NO";
    defparam add_33918_18.INJECT1_1 = "NO";
    CCU2D add_33918_16 (.A0(spi_byte_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48409), .COUT(n48410));
    defparam add_33918_16.INIT0 = 16'h5555;
    defparam add_33918_16.INIT1 = 16'h5555;
    defparam add_33918_16.INJECT1_0 = "NO";
    defparam add_33918_16.INJECT1_1 = "NO";
    CCU2D add_33918_14 (.A0(spi_byte_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48408), .COUT(n48409));
    defparam add_33918_14.INIT0 = 16'h5555;
    defparam add_33918_14.INIT1 = 16'h5555;
    defparam add_33918_14.INJECT1_0 = "NO";
    defparam add_33918_14.INJECT1_1 = "NO";
    CCU2D add_33918_12 (.A0(spi_byte_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48407), .COUT(n48408));
    defparam add_33918_12.INIT0 = 16'h5555;
    defparam add_33918_12.INIT1 = 16'h5555;
    defparam add_33918_12.INJECT1_0 = "NO";
    defparam add_33918_12.INJECT1_1 = "NO";
    CCU2D add_33918_10 (.A0(spi_byte_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48406), .COUT(n48407));
    defparam add_33918_10.INIT0 = 16'h5555;
    defparam add_33918_10.INIT1 = 16'h5555;
    defparam add_33918_10.INJECT1_0 = "NO";
    defparam add_33918_10.INJECT1_1 = "NO";
    CCU2D add_33918_8 (.A0(spi_byte_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48405), .COUT(n48406));
    defparam add_33918_8.INIT0 = 16'h5555;
    defparam add_33918_8.INIT1 = 16'h5555;
    defparam add_33918_8.INJECT1_0 = "NO";
    defparam add_33918_8.INJECT1_1 = "NO";
    CCU2D add_33918_6 (.A0(spi_byte_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48404), .COUT(n48405));
    defparam add_33918_6.INIT0 = 16'h5555;
    defparam add_33918_6.INIT1 = 16'h5555;
    defparam add_33918_6.INJECT1_0 = "NO";
    defparam add_33918_6.INJECT1_1 = "NO";
    CCU2D add_33918_4 (.A0(spi_byte_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48403), .COUT(n48404));
    defparam add_33918_4.INIT0 = 16'h5555;
    defparam add_33918_4.INIT1 = 16'h5555;
    defparam add_33918_4.INJECT1_0 = "NO";
    defparam add_33918_4.INJECT1_1 = "NO";
    CCU2D add_33918_2 (.A0(spi_byte_counter[1]), .B0(spi_byte_counter[0]), 
          .C0(GND_net), .D0(GND_net), .A1(spi_byte_counter[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n48403));
    defparam add_33918_2.INIT0 = 16'h7000;
    defparam add_33918_2.INIT1 = 16'h5555;
    defparam add_33918_2.INJECT1_0 = "NO";
    defparam add_33918_2.INJECT1_1 = "NO";
    LUT4 i24477_2_lut (.A(n55544), .B(n55545), .Z(n36657)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i24477_2_lut.init = 16'h8888;
    LUT4 i28797_2_lut (.A(delay_counter_31__N_659[2]), .B(n55544), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i28797_2_lut.init = 16'hbbbb;
    CCU2D add_33904_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48833), 
          .S0(n14501));
    defparam add_33904_cout.INIT0 = 16'h0000;
    defparam add_33904_cout.INIT1 = 16'h0000;
    defparam add_33904_cout.INJECT1_0 = "NO";
    defparam add_33904_cout.INJECT1_1 = "NO";
    CCU2D add_33904_31 (.A0(spi_byte_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48832), .COUT(n48833));
    defparam add_33904_31.INIT0 = 16'hf555;
    defparam add_33904_31.INIT1 = 16'h5555;
    defparam add_33904_31.INJECT1_0 = "NO";
    defparam add_33904_31.INJECT1_1 = "NO";
    CCU2D add_33904_29 (.A0(spi_byte_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48831), .COUT(n48832));
    defparam add_33904_29.INIT0 = 16'hf555;
    defparam add_33904_29.INIT1 = 16'hf555;
    defparam add_33904_29.INJECT1_0 = "NO";
    defparam add_33904_29.INJECT1_1 = "NO";
    CCU2D add_33904_27 (.A0(spi_byte_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48830), .COUT(n48831));
    defparam add_33904_27.INIT0 = 16'hf555;
    defparam add_33904_27.INIT1 = 16'hf555;
    defparam add_33904_27.INJECT1_0 = "NO";
    defparam add_33904_27.INJECT1_1 = "NO";
    CCU2D add_33904_25 (.A0(spi_byte_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48829), .COUT(n48830));
    defparam add_33904_25.INIT0 = 16'hf555;
    defparam add_33904_25.INIT1 = 16'hf555;
    defparam add_33904_25.INJECT1_0 = "NO";
    defparam add_33904_25.INJECT1_1 = "NO";
    LUT4 i2_4_lut_4_lut (.A(index[1]), .B(index[2]), .C(index[0]), .D(index[3]), 
         .Z(n50674)) /* synthesis lut_function=(!(A+(B (C+(D))+!B ((D)+!C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i2_4_lut_4_lut.init = 16'h0014;
    CCU2D add_33904_23 (.A0(spi_byte_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48828), .COUT(n48829));
    defparam add_33904_23.INIT0 = 16'hf555;
    defparam add_33904_23.INIT1 = 16'hf555;
    defparam add_33904_23.INJECT1_0 = "NO";
    defparam add_33904_23.INJECT1_1 = "NO";
    CCU2D add_33904_21 (.A0(spi_byte_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48827), .COUT(n48828));
    defparam add_33904_21.INIT0 = 16'hf555;
    defparam add_33904_21.INIT1 = 16'hf555;
    defparam add_33904_21.INJECT1_0 = "NO";
    defparam add_33904_21.INJECT1_1 = "NO";
    CCU2D add_33904_19 (.A0(spi_byte_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48826), .COUT(n48827));
    defparam add_33904_19.INIT0 = 16'hf555;
    defparam add_33904_19.INIT1 = 16'hf555;
    defparam add_33904_19.INJECT1_0 = "NO";
    defparam add_33904_19.INJECT1_1 = "NO";
    CCU2D add_33904_17 (.A0(spi_byte_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48825), .COUT(n48826));
    defparam add_33904_17.INIT0 = 16'hf555;
    defparam add_33904_17.INIT1 = 16'hf555;
    defparam add_33904_17.INJECT1_0 = "NO";
    defparam add_33904_17.INJECT1_1 = "NO";
    CCU2D add_33904_15 (.A0(spi_byte_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48824), .COUT(n48825));
    defparam add_33904_15.INIT0 = 16'hf555;
    defparam add_33904_15.INIT1 = 16'hf555;
    defparam add_33904_15.INJECT1_0 = "NO";
    defparam add_33904_15.INJECT1_1 = "NO";
    CCU2D add_33904_13 (.A0(spi_byte_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48823), .COUT(n48824));
    defparam add_33904_13.INIT0 = 16'hf555;
    defparam add_33904_13.INIT1 = 16'hf555;
    defparam add_33904_13.INJECT1_0 = "NO";
    defparam add_33904_13.INJECT1_1 = "NO";
    CCU2D add_33904_11 (.A0(spi_byte_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48822), .COUT(n48823));
    defparam add_33904_11.INIT0 = 16'hf555;
    defparam add_33904_11.INIT1 = 16'hf555;
    defparam add_33904_11.INJECT1_0 = "NO";
    defparam add_33904_11.INJECT1_1 = "NO";
    LUT4 mux_132_i4_3_lut (.A(index[3]), .B(DATA_OUT[4]), .C(n14326), 
         .Z(fb_31__N_715[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_132_i4_3_lut.init = 16'hcaca;
    CCU2D add_33904_9 (.A0(spi_byte_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48821), .COUT(n48822));
    defparam add_33904_9.INIT0 = 16'hf555;
    defparam add_33904_9.INIT1 = 16'hf555;
    defparam add_33904_9.INJECT1_0 = "NO";
    defparam add_33904_9.INJECT1_1 = "NO";
    CCU2D add_33904_7 (.A0(spi_byte_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48820), .COUT(n48821));
    defparam add_33904_7.INIT0 = 16'hf555;
    defparam add_33904_7.INIT1 = 16'hf555;
    defparam add_33904_7.INJECT1_0 = "NO";
    defparam add_33904_7.INJECT1_1 = "NO";
    CCU2D add_33904_5 (.A0(spi_byte_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48819), .COUT(n48820));
    defparam add_33904_5.INIT0 = 16'hf555;
    defparam add_33904_5.INIT1 = 16'hf555;
    defparam add_33904_5.INJECT1_0 = "NO";
    defparam add_33904_5.INJECT1_1 = "NO";
    CCU2D add_33904_3 (.A0(spi_byte_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_byte_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48818), .COUT(n48819));
    defparam add_33904_3.INIT0 = 16'hf555;
    defparam add_33904_3.INIT1 = 16'hf555;
    defparam add_33904_3.INJECT1_0 = "NO";
    defparam add_33904_3.INJECT1_1 = "NO";
    CCU2D add_33904_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(spi_byte_counter[0]), .B1(spi_byte_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48818));
    defparam add_33904_1.INIT0 = 16'hF000;
    defparam add_33904_1.INIT1 = 16'ha666;
    defparam add_33904_1.INJECT1_0 = "NO";
    defparam add_33904_1.INJECT1_1 = "NO";
    LUT4 mux_132_i3_3_lut (.A(index[2]), .B(DATA_OUT[3]), .C(n14326), 
         .Z(fb_31__N_715[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_132_i3_3_lut.init = 16'hcaca;
    LUT4 i28663_2_lut (.A(delay_counter_31__N_659[0]), .B(n55544), .Z(n1_adj_922)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(47[3] 113[12])
    defparam i28663_2_lut.init = 16'hbbbb;
    LUT4 mux_132_i2_3_lut (.A(index[1]), .B(DATA_OUT[2]), .C(n14326), 
         .Z(fb_31__N_715[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_132_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n54622), .B(n54681), .C(n54741), .D(n14431), .Z(sclk_c_enable_1283)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(31[12:17])
    defparam i1_4_lut.init = 16'h33b3;
    LUT4 mux_129_i1_3_lut (.A(n2[7]), .B(DATA_OUT[0]), .C(n14326), .Z(WrData_23__N_691[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_129_i1_3_lut.init = 16'hcaca;
    LUT4 i38619_4_lut (.A(n55545), .B(n7), .C(n14571), .D(n55544), .Z(sclk_c_enable_2505)) /* synthesis lut_function=(A+(B (C (D))+!B (C+!(D)))) */ ;
    defparam i38619_4_lut.init = 16'hfabb;
    LUT4 i1_2_lut_adj_882 (.A(n14326), .B(n14536), .Z(n7)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_882.init = 16'h8888;
    LUT4 i25019_1_lut (.A(n55544), .Z(n1_adj_923)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i25019_1_lut.init = 16'h5555;
    LUT4 i3_4_lut_adj_883 (.A(n54741), .B(spi_byte_counter[1]), .C(spi_byte_counter[2]), 
         .D(n131), .Z(n51592)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i3_4_lut_adj_883.init = 16'h2000;
    LUT4 mux_132_i1_3_lut (.A(index[0]), .B(DATA_OUT[1]), .C(n14326), 
         .Z(fb_31__N_715[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(53[5] 86[12])
    defparam mux_132_i1_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut (.A(index[0]), .B(index[1]), .C(index[3]), .D(index[2]), 
         .Z(n50606)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(54[24:29])
    defparam i3_3_lut_4_lut.init = 16'h0004;
    PFUMX i38975 (.BLUT(n55002), .ALUT(n55003), .C0(RX_RDY), .Z(sclk_c_enable_224));
    CCU2D add_3144_33 (.A0(delay_counter[31]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47834), .S0(delay_counter_31__N_659[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_33.INIT0 = 16'h5999;
    defparam add_3144_33.INIT1 = 16'h0000;
    defparam add_3144_33.INJECT1_0 = "NO";
    defparam add_3144_33.INJECT1_1 = "NO";
    CCU2D add_3144_31 (.A0(delay_counter[29]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47833), .COUT(n47834), .S0(delay_counter_31__N_659[29]), 
          .S1(delay_counter_31__N_659[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_31.INIT0 = 16'h5999;
    defparam add_3144_31.INIT1 = 16'h5999;
    defparam add_3144_31.INJECT1_0 = "NO";
    defparam add_3144_31.INJECT1_1 = "NO";
    CCU2D add_3144_29 (.A0(delay_counter[27]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47832), .COUT(n47833), .S0(delay_counter_31__N_659[27]), 
          .S1(delay_counter_31__N_659[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_29.INIT0 = 16'h5999;
    defparam add_3144_29.INIT1 = 16'h5999;
    defparam add_3144_29.INJECT1_0 = "NO";
    defparam add_3144_29.INJECT1_1 = "NO";
    CCU2D add_3144_27 (.A0(delay_counter[25]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47831), .COUT(n47832), .S0(delay_counter_31__N_659[25]), 
          .S1(delay_counter_31__N_659[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_27.INIT0 = 16'h5999;
    defparam add_3144_27.INIT1 = 16'h5999;
    defparam add_3144_27.INJECT1_0 = "NO";
    defparam add_3144_27.INJECT1_1 = "NO";
    CCU2D add_3144_25 (.A0(delay_counter[23]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47830), .COUT(n47831), .S0(delay_counter_31__N_659[23]), 
          .S1(delay_counter_31__N_659[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_25.INIT0 = 16'h5999;
    defparam add_3144_25.INIT1 = 16'h5999;
    defparam add_3144_25.INJECT1_0 = "NO";
    defparam add_3144_25.INJECT1_1 = "NO";
    CCU2D add_3144_23 (.A0(delay_counter[21]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47829), .COUT(n47830), .S0(delay_counter_31__N_659[21]), 
          .S1(delay_counter_31__N_659[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_23.INIT0 = 16'h5999;
    defparam add_3144_23.INIT1 = 16'h5999;
    defparam add_3144_23.INJECT1_0 = "NO";
    defparam add_3144_23.INJECT1_1 = "NO";
    CCU2D add_3144_21 (.A0(delay_counter[19]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47828), .COUT(n47829), .S0(delay_counter_31__N_659[19]), 
          .S1(delay_counter_31__N_659[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_21.INIT0 = 16'h5999;
    defparam add_3144_21.INIT1 = 16'h5999;
    defparam add_3144_21.INJECT1_0 = "NO";
    defparam add_3144_21.INJECT1_1 = "NO";
    CCU2D add_3144_19 (.A0(delay_counter[17]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47827), .COUT(n47828), .S0(delay_counter_31__N_659[17]), 
          .S1(delay_counter_31__N_659[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_19.INIT0 = 16'h5999;
    defparam add_3144_19.INIT1 = 16'h5999;
    defparam add_3144_19.INJECT1_0 = "NO";
    defparam add_3144_19.INJECT1_1 = "NO";
    CCU2D add_3144_17 (.A0(delay_counter[15]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47826), .COUT(n47827), .S0(delay_counter_31__N_659[15]), 
          .S1(delay_counter_31__N_659[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_17.INIT0 = 16'h5999;
    defparam add_3144_17.INIT1 = 16'h5999;
    defparam add_3144_17.INJECT1_0 = "NO";
    defparam add_3144_17.INJECT1_1 = "NO";
    CCU2D add_3144_15 (.A0(delay_counter[13]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47825), .COUT(n47826), .S0(delay_counter_31__N_659[13]), 
          .S1(delay_counter_31__N_659[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_15.INIT0 = 16'h5999;
    defparam add_3144_15.INIT1 = 16'h5999;
    defparam add_3144_15.INJECT1_0 = "NO";
    defparam add_3144_15.INJECT1_1 = "NO";
    CCU2D add_3144_13 (.A0(delay_counter[11]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47824), .COUT(n47825), .S0(delay_counter_31__N_659[11]), 
          .S1(delay_counter_31__N_659[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_13.INIT0 = 16'h5999;
    defparam add_3144_13.INIT1 = 16'h5999;
    defparam add_3144_13.INJECT1_0 = "NO";
    defparam add_3144_13.INJECT1_1 = "NO";
    CCU2D add_3144_11 (.A0(delay_counter[9]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47823), .COUT(n47824), .S0(delay_counter_31__N_659[9]), 
          .S1(delay_counter_31__N_659[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_11.INIT0 = 16'h5999;
    defparam add_3144_11.INIT1 = 16'h5999;
    defparam add_3144_11.INJECT1_0 = "NO";
    defparam add_3144_11.INJECT1_1 = "NO";
    CCU2D add_3144_9 (.A0(delay_counter[7]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47822), .COUT(n47823), .S0(delay_counter_31__N_659[7]), 
          .S1(delay_counter_31__N_659[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_9.INIT0 = 16'h5999;
    defparam add_3144_9.INIT1 = 16'h5999;
    defparam add_3144_9.INJECT1_0 = "NO";
    defparam add_3144_9.INJECT1_1 = "NO";
    CCU2D add_3144_7 (.A0(delay_counter[5]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47821), .COUT(n47822), .S0(delay_counter_31__N_659[5]), 
          .S1(delay_counter_31__N_659[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_7.INIT0 = 16'h5999;
    defparam add_3144_7.INIT1 = 16'h5999;
    defparam add_3144_7.INJECT1_0 = "NO";
    defparam add_3144_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_884 (.A(n55545), .B(n14326), .C(RX_RDY), .Z(SPI_CS_N_880)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam i1_3_lut_adj_884.init = 16'h5151;
    CCU2D add_3144_5 (.A0(delay_counter[3]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47820), .COUT(n47821), .S0(delay_counter_31__N_659[3]), 
          .S1(delay_counter_31__N_659[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_5.INIT0 = 16'h5999;
    defparam add_3144_5.INIT1 = 16'h5999;
    defparam add_3144_5.INJECT1_0 = "NO";
    defparam add_3144_5.INJECT1_1 = "NO";
    CCU2D add_3144_3 (.A0(delay_counter[1]), .B0(n14571), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(n14571), .C1(GND_net), 
          .D1(GND_net), .CIN(n47819), .COUT(n47820), .S0(delay_counter_31__N_659[1]), 
          .S1(delay_counter_31__N_659[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_3.INIT0 = 16'h5999;
    defparam add_3144_3.INIT1 = 16'h5999;
    defparam add_3144_3.INJECT1_0 = "NO";
    defparam add_3144_3.INJECT1_1 = "NO";
    CCU2D add_3144_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(n14571), .C1(GND_net), .D1(GND_net), 
          .COUT(n47819), .S1(delay_counter_31__N_659[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(97[5] 102[12])
    defparam add_3144_1.INIT0 = 16'hF000;
    defparam add_3144_1.INIT1 = 16'h5999;
    defparam add_3144_1.INJECT1_0 = "NO";
    defparam add_3144_1.INJECT1_1 = "NO";
    FD1P3IX state_i1_rep_850 (.D(state[0]), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(sclk_c_enable_1092)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i1_rep_850.GSR = "DISABLED";
    FD1P3IX state_i1_rep_848 (.D(state[0]), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(n55547)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i1_rep_848.GSR = "DISABLED";
    FD1P3IX state_i1_rep_847 (.D(state[0]), .SP(sclk_c_enable_2505), .CD(state[1]), 
            .CK(sclk_c), .Q(sclk_c_enable_1028)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i1_rep_847.GSR = "DISABLED";
    FD1P3IX state_i1_rep_846 (.D(state[0]), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1092), 
            .CK(sclk_c), .Q(n55545)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i1_rep_846.GSR = "DISABLED";
    FD1P3IX state_i0_rep_845 (.D(n1_adj_923), .SP(sclk_c_enable_2505), .CD(sclk_c_enable_1028), 
            .CK(sclk_c), .Q(n55544)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=14, LSE_RCOL=22, LSE_LLINE=359, LSE_RLINE=359 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/load_mem.vhd(29[2] 114[14])
    defparam state_i0_rep_845.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U30 
//

module \WS2812(48000000,"111111111")_U30  (sclk_c, \port_status[18] , ws2813_out_c_18, 
            \Q[18] , \RdAddress[18] , GND_net);
    input sclk_c;
    output \port_status[18] ;
    output ws2813_out_c_18;
    input [23:0]\Q[18] ;
    output [8:0]\RdAddress[18] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1650;
    wire [31:0]n10660;
    
    wire sclk_c_enable_162, n54753, sclk_c_enable_163, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_166;
    wire [2:0]state_2__N_104;
    
    wire n14151, n6909, n53199, n53200;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53203;
    wire [31:0]n447;
    
    wire n54972, n54971, n53201, n53202, n53204, n53205, n53368, 
        serial_N_437, n53366, n53367;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1468, n36448;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1435;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1499;
    wire [31:0]bit_counter_31__N_172;
    
    wire n54561, n54767, n54699;
    wire [31:0]n10484;
    
    wire n54690, n14116, n76, n42688;
    wire [8:0]n118;
    
    wire n53364, n53365, n68;
    wire [6:0]n15121;
    
    wire n10659, n52679, n37607, n4, n54572, n54634, n103, n53362, 
        n53191, n53192, n53193, n53194, n1, n1_adj_915, n53195, 
        n53196, n53197, n53198, n54632, n54887, n36266, n54886, 
        n54888, n36270, n53363, n54973;
    wire [31:0]bit_counter_31__N_204;
    
    wire n47898, n47897, n47896, n47895, n47894, n47893, n47892, 
        n69, n47891, n47890, n47889, n47888, n47887, n47886, n47885, 
        n47884, n47883, n15, n14, n48104, n48103, n48102, n48101, 
        n48100, n48099, n48817, n48816, n48815, n48814, n48813, 
        n48812, n48811, n48810, n48809, n48808, n48807, n48806, 
        n48805, n48804, n48803, n48802, n48098, n48097, n48096, 
        n48095, n48094, n48093, n48092, n48091, n48090, n48089, 
        n48087, n48086, n48085, n48084, n48769, n48768, n48767, 
        n48766, n48765, n48764, n48763, n48762, n48761, n48760, 
        n48759, n48758, n48757, n48756, n48755, n48754;
    
    FD1P3AX delay_counter_i0_i0 (.D(n10660[0]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54753), .SP(sclk_c_enable_162), .CK(sclk_c), 
            .Q(\port_status[18] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_163), .CK(sclk_c), 
            .Q(ws2813_out_c_18)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_166), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_166), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_166), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n14151), .Z(n6909)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 i38458_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n14151), .Z(sclk_c_enable_166)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38458_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    L6MUX21 i37997 (.D0(n53199), .D1(n53200), .SD(bit_counter[2]), .Z(n53203));
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 mux_2894_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n14151), .Z(n54972)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2894_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2894_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n14151), .Z(n54971)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2894_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    L6MUX21 i37998 (.D0(n53201), .D1(n53202), .SD(bit_counter[2]), .Z(n53204));
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53205), .B(n53368), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    L6MUX21 i38162 (.D0(n53366), .D1(n53367), .SD(bit_counter[2]), .Z(n53368));
    FD1P3IX pixel_i0 (.D(\Q[18] [0]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n54561), .B(n54767), .C(n447[7]), .D(n54699), 
         .Z(n10484[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_799 (.A(n54561), .B(n54767), .C(n447[8]), 
         .D(n54699), .Z(n10484[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_799.init = 16'hf888;
    LUT4 mux_2083_i2_4_lut_4_lut (.A(n54690), .B(n54699), .C(n6909), .D(n14116), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2083_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 i1_3_lut_4_lut_adj_800 (.A(n54561), .B(n54767), .C(n447[9]), 
         .D(n54699), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_800.init = 16'hf888;
    FD1P3AX delay_counter_i0_i1 (.D(n10660[1]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n10660[3]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n10660[7]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n10660[8]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n10660[9]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n10660[12]), .SP(sclk_c_enable_1650), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n42688), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_801 (.A(state[2]), .B(n42688), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_801.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_802 (.A(state[2]), .B(n42688), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_802.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_803 (.A(state[2]), .B(n42688), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_803.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_804 (.A(state[2]), .B(n42688), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_804.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_805 (.A(state[2]), .B(n42688), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_805.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_806 (.A(state[2]), .B(n42688), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_806.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_807 (.A(state[2]), .B(n42688), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_807.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_808 (.A(state[2]), .B(n42688), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_808.init = 16'h1010;
    PFUMX i38161 (.BLUT(n53364), .ALUT(n53365), .C0(bit_counter[1]), .Z(n53367));
    LUT4 mux_2904_i2_4_lut (.A(n68), .B(n15121[0]), .C(n10659), .D(n52679), 
         .Z(n10660[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2904_i4_4_lut (.A(n37607), .B(n54690), .C(n10659), .D(n4), 
         .Z(n10660[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42688), .B(n54572), .C(n447[3]), .D(n54699), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2904_i8_4_lut (.A(n10484[7]), .B(n54690), .C(n10659), .D(n54572), 
         .Z(n10660[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i8_4_lut.init = 16'h303a;
    LUT4 mux_2083_i1_4_lut (.A(n54634), .B(n54690), .C(n6909), .D(n54699), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2083_i1_4_lut.init = 16'h3f3a;
    LUT4 mux_2904_i9_4_lut (.A(n10484[8]), .B(n54690), .C(n10659), .D(n54572), 
         .Z(n10660[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i9_4_lut.init = 16'h303a;
    FD1P3IX pixel_i23 (.D(\Q[18] [23]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[18] [22]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[18] [21]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[18] [20]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[18] [19]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[18] [18]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[18] [17]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[18] [16]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[18] [15]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[18] [14]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[18] [13]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[18] [12]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[18] [11]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[18] [10]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[18] [9]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[18] [8]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[18] [7]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[18] [6]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[18] [5]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[18] [4]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[18] [3]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[18] [2]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[18] [1]), .SP(sclk_c_enable_1468), .CD(n36448), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1435), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54634), .C(n14151), .D(n54767), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    LUT4 mux_2904_i10_4_lut (.A(n76), .B(n54690), .C(n10659), .D(n54572), 
         .Z(n10660[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i10_4_lut.init = 16'h303a;
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    LUT4 mux_2904_i13_4_lut (.A(n54572), .B(n54690), .C(n10659), .D(n103), 
         .Z(n10660[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i13_4_lut.init = 16'h3530;
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1468), 
            .CD(n36448), .CK(sclk_c), .Q(\RdAddress[18] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    LUT4 i38156_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38156_3_lut.init = 16'hcaca;
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    PFUMX i37993 (.BLUT(n53191), .ALUT(n53192), .C0(bit_counter[1]), .Z(n53199));
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    PFUMX i37994 (.BLUT(n53193), .ALUT(n53194), .C0(bit_counter[1]), .Z(n53200));
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1499), .CD(n36448), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_915), .SP(sclk_c_enable_1499), .CD(n36448), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    PFUMX i37995 (.BLUT(n53195), .ALUT(n53196), .C0(bit_counter[1]), .Z(n53201));
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1499), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    PFUMX i37996 (.BLUT(n53197), .ALUT(n53198), .C0(bit_counter[1]), .Z(n53202));
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54767), .B(state[1]), .C(n54634), .D(n54632), 
         .Z(n52679)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 mux_2894_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14151), .Z(n54887)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2894_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 i24054_2_lut_4_lut (.A(n54632), .B(state[0]), .C(state[1]), .D(n10659), 
         .Z(n36266)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i24054_2_lut_4_lut.init = 16'hfd00;
    LUT4 mux_2894_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14116), .Z(n54886)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2894_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i37992_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37992_3_lut.init = 16'hcaca;
    LUT4 i37991_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37991_3_lut.init = 16'hcaca;
    LUT4 i37990_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37990_3_lut.init = 16'hcaca;
    LUT4 i37989_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37989_3_lut.init = 16'hcaca;
    LUT4 i37988_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37988_3_lut.init = 16'hcaca;
    LUT4 i37987_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37987_3_lut.init = 16'hcaca;
    LUT4 i37986_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37986_3_lut.init = 16'hcaca;
    LUT4 i37985_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37985_3_lut.init = 16'hcaca;
    PFUMX i38899 (.BLUT(n54886), .ALUT(n54887), .C0(state[1]), .Z(n54888));
    L6MUX21 i37999 (.D0(n53203), .D1(n53204), .SD(bit_counter[3]), .Z(n53205));
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    PFUMX i38160 (.BLUT(n53362), .ALUT(n53363), .C0(bit_counter[1]), .Z(n53366));
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1650), 
            .CD(n36270), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1650), .CD(n36270), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1650), .CD(n36270), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54973), .SP(sclk_c_enable_1650), .CD(n36266), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54888), .SP(sclk_c_enable_1650), .CD(n36266), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=333, LSE_RLINE=333 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i38159_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38159_3_lut.init = 16'hcaca;
    LUT4 i38158_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38158_3_lut.init = 16'hcaca;
    LUT4 i38157_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38157_3_lut.init = 16'hcaca;
    LUT4 i38428_2_lut_rep_749 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1499)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38428_2_lut_rep_749.init = 16'h9999;
    LUT4 i25402_1_lut_rep_750 (.A(state[2]), .Z(n54753)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25402_1_lut_rep_750.init = 16'h5555;
    LUT4 i29965_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i29965_3_lut_3_lut.init = 16'h5151;
    LUT4 i28792_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28792_2_lut.init = 16'hbbbb;
    LUT4 i28791_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_915)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28791_2_lut.init = 16'hbbbb;
    CCU2D add_3138_33 (.A0(bit_counter[31]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47898), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_33.INIT0 = 16'h5999;
    defparam add_3138_33.INIT1 = 16'h0000;
    defparam add_3138_33.INJECT1_0 = "NO";
    defparam add_3138_33.INJECT1_1 = "NO";
    CCU2D add_3138_31 (.A0(bit_counter[29]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47897), .COUT(n47898), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_31.INIT0 = 16'h5999;
    defparam add_3138_31.INIT1 = 16'h5999;
    defparam add_3138_31.INJECT1_0 = "NO";
    defparam add_3138_31.INJECT1_1 = "NO";
    CCU2D add_3138_29 (.A0(bit_counter[27]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47896), .COUT(n47897), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_29.INIT0 = 16'h5999;
    defparam add_3138_29.INIT1 = 16'h5999;
    defparam add_3138_29.INJECT1_0 = "NO";
    defparam add_3138_29.INJECT1_1 = "NO";
    CCU2D add_3138_27 (.A0(bit_counter[25]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47895), .COUT(n47896), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_27.INIT0 = 16'h5999;
    defparam add_3138_27.INIT1 = 16'h5999;
    defparam add_3138_27.INJECT1_0 = "NO";
    defparam add_3138_27.INJECT1_1 = "NO";
    CCU2D add_3138_25 (.A0(bit_counter[23]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47894), .COUT(n47895), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_25.INIT0 = 16'h5999;
    defparam add_3138_25.INIT1 = 16'h5999;
    defparam add_3138_25.INJECT1_0 = "NO";
    defparam add_3138_25.INJECT1_1 = "NO";
    CCU2D add_3138_23 (.A0(bit_counter[21]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47893), .COUT(n47894), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_23.INIT0 = 16'h5999;
    defparam add_3138_23.INIT1 = 16'h5999;
    defparam add_3138_23.INJECT1_0 = "NO";
    defparam add_3138_23.INJECT1_1 = "NO";
    CCU2D add_3138_21 (.A0(bit_counter[19]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47892), .COUT(n47893), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_21.INIT0 = 16'h5999;
    defparam add_3138_21.INIT1 = 16'h5999;
    defparam add_3138_21.INJECT1_0 = "NO";
    defparam add_3138_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_696_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54699)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_696_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_809 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_809.init = 16'he0f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n14151), 
         .Z(sclk_c_enable_163)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_rep_687_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54690)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_687_3_lut.init = 16'hf8f8;
    CCU2D add_3138_19 (.A0(bit_counter[17]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47891), .COUT(n47892), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_19.INIT0 = 16'h5999;
    defparam add_3138_19.INIT1 = 16'h5999;
    defparam add_3138_19.INJECT1_0 = "NO";
    defparam add_3138_19.INJECT1_1 = "NO";
    CCU2D add_3138_17 (.A0(bit_counter[15]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47890), .COUT(n47891), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_17.INIT0 = 16'h5999;
    defparam add_3138_17.INIT1 = 16'h5999;
    defparam add_3138_17.INJECT1_0 = "NO";
    defparam add_3138_17.INJECT1_1 = "NO";
    LUT4 i24299_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36448)) /* synthesis lut_function=(A (B)) */ ;
    defparam i24299_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    CCU2D add_3138_15 (.A0(bit_counter[13]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47889), .COUT(n47890), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_15.INIT0 = 16'h5999;
    defparam add_3138_15.INIT1 = 16'h5999;
    defparam add_3138_15.INJECT1_0 = "NO";
    defparam add_3138_15.INJECT1_1 = "NO";
    LUT4 i24078_4_lut (.A(sclk_c_enable_1650), .B(n54699), .C(n10659), 
         .D(n54572), .Z(n36270)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i24078_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_adj_810 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15121[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_810.init = 16'h7070;
    LUT4 i1_3_lut_rep_689_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1468)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_689_4_lut_3_lut.init = 16'h8989;
    CCU2D add_3138_13 (.A0(bit_counter[11]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47888), .COUT(n47889), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_13.INIT0 = 16'h5999;
    defparam add_3138_13.INIT1 = 16'h5999;
    defparam add_3138_13.INJECT1_0 = "NO";
    defparam add_3138_13.INJECT1_1 = "NO";
    CCU2D add_3138_11 (.A0(bit_counter[9]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47887), .COUT(n47888), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_11.INIT0 = 16'h5999;
    defparam add_3138_11.INIT1 = 16'h5999;
    defparam add_3138_11.INJECT1_0 = "NO";
    defparam add_3138_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_764 (.A(state[0]), .B(state[2]), .Z(n54767)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_764.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_811 (.A(state[0]), .B(state[2]), .C(n14116), 
         .D(state[1]), .Z(n37607)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_811.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n14116), 
         .D(state[1]), .Z(sclk_c_enable_1435)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_812 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_812.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_813 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_813.init = 16'h2020;
    CCU2D add_3138_9 (.A0(bit_counter[7]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47886), .COUT(n47887), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_9.INIT0 = 16'h5999;
    defparam add_3138_9.INIT1 = 16'h5999;
    defparam add_3138_9.INJECT1_0 = "NO";
    defparam add_3138_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_814 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_814.init = 16'h2020;
    CCU2D add_3138_7 (.A0(bit_counter[5]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47885), .COUT(n47886), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_7.INIT0 = 16'h5999;
    defparam add_3138_7.INIT1 = 16'h5999;
    defparam add_3138_7.INJECT1_0 = "NO";
    defparam add_3138_7.INJECT1_1 = "NO";
    CCU2D add_3138_5 (.A0(bit_counter[3]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47884), .COUT(n47885), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_5.INIT0 = 16'h5999;
    defparam add_3138_5.INIT1 = 16'h5999;
    defparam add_3138_5.INJECT1_0 = "NO";
    defparam add_3138_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_815 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_815.init = 16'h2020;
    CCU2D add_3138_3 (.A0(bit_counter[1]), .B0(n14116), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n14116), .C1(GND_net), 
          .D1(GND_net), .CIN(n47883), .COUT(n47884), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_3.INIT0 = 16'h5999;
    defparam add_3138_3.INIT1 = 16'h5999;
    defparam add_3138_3.INJECT1_0 = "NO";
    defparam add_3138_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_816 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_816.init = 16'h2020;
    CCU2D add_3138_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n14116), .C1(GND_net), .D1(GND_net), 
          .COUT(n47883), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3138_1.INIT0 = 16'hF000;
    defparam add_3138_1.INIT1 = 16'h5999;
    defparam add_3138_1.INJECT1_0 = "NO";
    defparam add_3138_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_817 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_817.init = 16'h2020;
    LUT4 mux_2904_i1_4_lut (.A(n69), .B(n15121[0]), .C(n10659), .D(n52679), 
         .Z(n10660[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2904_i1_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_3_lut_adj_818 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_818.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_819 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_819.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_820 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_820.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_821 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_821.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_822 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_822.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_823 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_823.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_824 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_824.init = 16'h2020;
    LUT4 i2916_3_lut (.A(state[2]), .B(state[1]), .C(n14151), .Z(n10659)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2916_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_3_lut_adj_825 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_825.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_826 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_826.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_827 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_827.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_828 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_828.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_829 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_829.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_830 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_830.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_831 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_831.init = 16'h2020;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42688)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_832 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_832.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_833 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_833.init = 16'h2020;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_834 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_834.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_835 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_835.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_836 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_836.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_837 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_837.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_838 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_838.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_839 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_839.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_840 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_840.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_841 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_841.init = 16'h2020;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48104), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48103), .COUT(n48104), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48102), .COUT(n48103), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48101), .COUT(n48102), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48100), .COUT(n48101), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48099), .COUT(n48100), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_33936_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48817), 
          .S0(n14151));
    defparam add_33936_cout.INIT0 = 16'h0000;
    defparam add_33936_cout.INIT1 = 16'h0000;
    defparam add_33936_cout.INJECT1_0 = "NO";
    defparam add_33936_cout.INJECT1_1 = "NO";
    CCU2D add_33936_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48816), .COUT(n48817));
    defparam add_33936_31.INIT0 = 16'hf555;
    defparam add_33936_31.INIT1 = 16'h5555;
    defparam add_33936_31.INJECT1_0 = "NO";
    defparam add_33936_31.INJECT1_1 = "NO";
    CCU2D add_33936_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48815), .COUT(n48816));
    defparam add_33936_29.INIT0 = 16'hf555;
    defparam add_33936_29.INIT1 = 16'hf555;
    defparam add_33936_29.INJECT1_0 = "NO";
    defparam add_33936_29.INJECT1_1 = "NO";
    CCU2D add_33936_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48814), .COUT(n48815));
    defparam add_33936_27.INIT0 = 16'hf555;
    defparam add_33936_27.INIT1 = 16'hf555;
    defparam add_33936_27.INJECT1_0 = "NO";
    defparam add_33936_27.INJECT1_1 = "NO";
    CCU2D add_33936_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48813), .COUT(n48814));
    defparam add_33936_25.INIT0 = 16'hf555;
    defparam add_33936_25.INIT1 = 16'hf555;
    defparam add_33936_25.INJECT1_0 = "NO";
    defparam add_33936_25.INJECT1_1 = "NO";
    CCU2D add_33936_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48812), .COUT(n48813));
    defparam add_33936_23.INIT0 = 16'hf555;
    defparam add_33936_23.INIT1 = 16'hf555;
    defparam add_33936_23.INJECT1_0 = "NO";
    defparam add_33936_23.INJECT1_1 = "NO";
    CCU2D add_33936_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48811), .COUT(n48812));
    defparam add_33936_21.INIT0 = 16'hf555;
    defparam add_33936_21.INIT1 = 16'hf555;
    defparam add_33936_21.INJECT1_0 = "NO";
    defparam add_33936_21.INJECT1_1 = "NO";
    CCU2D add_33936_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48810), .COUT(n48811));
    defparam add_33936_19.INIT0 = 16'hf555;
    defparam add_33936_19.INIT1 = 16'hf555;
    defparam add_33936_19.INJECT1_0 = "NO";
    defparam add_33936_19.INJECT1_1 = "NO";
    CCU2D add_33936_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48809), .COUT(n48810));
    defparam add_33936_17.INIT0 = 16'hf555;
    defparam add_33936_17.INIT1 = 16'hf555;
    defparam add_33936_17.INJECT1_0 = "NO";
    defparam add_33936_17.INJECT1_1 = "NO";
    CCU2D add_33936_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48808), .COUT(n48809));
    defparam add_33936_15.INIT0 = 16'hf555;
    defparam add_33936_15.INIT1 = 16'hf555;
    defparam add_33936_15.INJECT1_0 = "NO";
    defparam add_33936_15.INJECT1_1 = "NO";
    CCU2D add_33936_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48807), .COUT(n48808));
    defparam add_33936_13.INIT0 = 16'hf555;
    defparam add_33936_13.INIT1 = 16'hf555;
    defparam add_33936_13.INJECT1_0 = "NO";
    defparam add_33936_13.INJECT1_1 = "NO";
    CCU2D add_33936_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48806), .COUT(n48807));
    defparam add_33936_11.INIT0 = 16'hf555;
    defparam add_33936_11.INIT1 = 16'hf555;
    defparam add_33936_11.INJECT1_0 = "NO";
    defparam add_33936_11.INJECT1_1 = "NO";
    CCU2D add_33936_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48805), .COUT(n48806));
    defparam add_33936_9.INIT0 = 16'hf555;
    defparam add_33936_9.INIT1 = 16'hf555;
    defparam add_33936_9.INJECT1_0 = "NO";
    defparam add_33936_9.INJECT1_1 = "NO";
    CCU2D add_33936_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48804), .COUT(n48805));
    defparam add_33936_7.INIT0 = 16'hf555;
    defparam add_33936_7.INIT1 = 16'hf555;
    defparam add_33936_7.INJECT1_0 = "NO";
    defparam add_33936_7.INJECT1_1 = "NO";
    CCU2D add_33936_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48803), .COUT(n48804));
    defparam add_33936_5.INIT0 = 16'hf555;
    defparam add_33936_5.INIT1 = 16'hf555;
    defparam add_33936_5.INJECT1_0 = "NO";
    defparam add_33936_5.INJECT1_1 = "NO";
    CCU2D add_33936_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48802), .COUT(n48803));
    defparam add_33936_3.INIT0 = 16'hf555;
    defparam add_33936_3.INIT1 = 16'hf555;
    defparam add_33936_3.INJECT1_0 = "NO";
    defparam add_33936_3.INJECT1_1 = "NO";
    CCU2D add_33936_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48802));
    defparam add_33936_1.INIT0 = 16'hF000;
    defparam add_33936_1.INIT1 = 16'ha666;
    defparam add_33936_1.INJECT1_0 = "NO";
    defparam add_33936_1.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48098), .COUT(n48099), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48097), .COUT(n48098), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48096), .COUT(n48097), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48095), .COUT(n48096), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48094), .COUT(n48095), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48093), .COUT(n48094), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48092), .COUT(n48093), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48091), .COUT(n48092), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48090), .COUT(n48091), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48089), .COUT(n48090), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48089), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48087), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48086), .COUT(n48087), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48085), .COUT(n48086), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48084), .COUT(n48085), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48084), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_33938_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48769), 
          .S0(n14116));
    defparam add_33938_cout.INIT0 = 16'h0000;
    defparam add_33938_cout.INIT1 = 16'h0000;
    defparam add_33938_cout.INJECT1_0 = "NO";
    defparam add_33938_cout.INJECT1_1 = "NO";
    CCU2D add_33938_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48768), .COUT(n48769));
    defparam add_33938_31.INIT0 = 16'hf555;
    defparam add_33938_31.INIT1 = 16'h5555;
    defparam add_33938_31.INJECT1_0 = "NO";
    defparam add_33938_31.INJECT1_1 = "NO";
    CCU2D add_33938_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48767), .COUT(n48768));
    defparam add_33938_29.INIT0 = 16'hf555;
    defparam add_33938_29.INIT1 = 16'hf555;
    defparam add_33938_29.INJECT1_0 = "NO";
    defparam add_33938_29.INJECT1_1 = "NO";
    CCU2D add_33938_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48766), .COUT(n48767));
    defparam add_33938_27.INIT0 = 16'hf555;
    defparam add_33938_27.INIT1 = 16'hf555;
    defparam add_33938_27.INJECT1_0 = "NO";
    defparam add_33938_27.INJECT1_1 = "NO";
    CCU2D add_33938_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48765), .COUT(n48766));
    defparam add_33938_25.INIT0 = 16'hf555;
    defparam add_33938_25.INIT1 = 16'hf555;
    defparam add_33938_25.INJECT1_0 = "NO";
    defparam add_33938_25.INJECT1_1 = "NO";
    CCU2D add_33938_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48764), .COUT(n48765));
    defparam add_33938_23.INIT0 = 16'hf555;
    defparam add_33938_23.INIT1 = 16'hf555;
    defparam add_33938_23.INJECT1_0 = "NO";
    defparam add_33938_23.INJECT1_1 = "NO";
    CCU2D add_33938_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48763), .COUT(n48764));
    defparam add_33938_21.INIT0 = 16'hf555;
    defparam add_33938_21.INIT1 = 16'hf555;
    defparam add_33938_21.INJECT1_0 = "NO";
    defparam add_33938_21.INJECT1_1 = "NO";
    CCU2D add_33938_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48762), .COUT(n48763));
    defparam add_33938_19.INIT0 = 16'hf555;
    defparam add_33938_19.INIT1 = 16'hf555;
    defparam add_33938_19.INJECT1_0 = "NO";
    defparam add_33938_19.INJECT1_1 = "NO";
    CCU2D add_33938_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48761), .COUT(n48762));
    defparam add_33938_17.INIT0 = 16'hf555;
    defparam add_33938_17.INIT1 = 16'hf555;
    defparam add_33938_17.INJECT1_0 = "NO";
    defparam add_33938_17.INJECT1_1 = "NO";
    CCU2D add_33938_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48760), .COUT(n48761));
    defparam add_33938_15.INIT0 = 16'hf555;
    defparam add_33938_15.INIT1 = 16'hf555;
    defparam add_33938_15.INJECT1_0 = "NO";
    defparam add_33938_15.INJECT1_1 = "NO";
    CCU2D add_33938_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48759), .COUT(n48760));
    defparam add_33938_13.INIT0 = 16'hf555;
    defparam add_33938_13.INIT1 = 16'hf555;
    defparam add_33938_13.INJECT1_0 = "NO";
    defparam add_33938_13.INJECT1_1 = "NO";
    CCU2D add_33938_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48758), .COUT(n48759));
    defparam add_33938_11.INIT0 = 16'hf555;
    defparam add_33938_11.INIT1 = 16'hf555;
    defparam add_33938_11.INJECT1_0 = "NO";
    defparam add_33938_11.INJECT1_1 = "NO";
    CCU2D add_33938_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48757), .COUT(n48758));
    defparam add_33938_9.INIT0 = 16'hf555;
    defparam add_33938_9.INIT1 = 16'hf555;
    defparam add_33938_9.INJECT1_0 = "NO";
    defparam add_33938_9.INJECT1_1 = "NO";
    CCU2D add_33938_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48756), .COUT(n48757));
    defparam add_33938_7.INIT0 = 16'hf555;
    defparam add_33938_7.INIT1 = 16'hf555;
    defparam add_33938_7.INJECT1_0 = "NO";
    defparam add_33938_7.INJECT1_1 = "NO";
    CCU2D add_33938_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48755), .COUT(n48756));
    defparam add_33938_5.INIT0 = 16'hf555;
    defparam add_33938_5.INIT1 = 16'hf555;
    defparam add_33938_5.INJECT1_0 = "NO";
    defparam add_33938_5.INJECT1_1 = "NO";
    CCU2D add_33938_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48754), .COUT(n48755));
    defparam add_33938_3.INIT0 = 16'hf555;
    defparam add_33938_3.INIT1 = 16'hf555;
    defparam add_33938_3.INJECT1_0 = "NO";
    defparam add_33938_3.INJECT1_1 = "NO";
    CCU2D add_33938_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48754));
    defparam add_33938_1.INIT0 = 16'hF000;
    defparam add_33938_1.INIT1 = 16'ha666;
    defparam add_33938_1.INJECT1_0 = "NO";
    defparam add_33938_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_629 (.A(state[2]), .B(n14151), .Z(n54632)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_629.init = 16'h4444;
    LUT4 i1_2_lut_rep_569_3_lut (.A(state[2]), .B(n14151), .C(state[1]), 
         .Z(n54572)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_569_3_lut.init = 16'h4040;
    LUT4 i107_3_lut_4_lut (.A(n42688), .B(n14116), .C(n54699), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 i38574_3_lut_rep_570_4_lut (.A(state[2]), .B(n14151), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1650)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38574_3_lut_rep_570_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_rep_631 (.A(n42688), .B(n14116), .Z(n54634)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_631.init = 16'h8888;
    PFUMX i38955 (.BLUT(n54971), .ALUT(n54972), .C0(state[0]), .Z(n54973));
    LUT4 i1_2_lut_rep_558_3_lut (.A(n42688), .B(n14116), .C(state[1]), 
         .Z(n54561)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_558_3_lut.init = 16'h0808;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \WS2812(48000000,"111111111")_U29 
//

module \WS2812(48000000,"111111111")_U29  (sclk_c, \port_status[19] , ws2813_out_c_19, 
            \Q[19] , \RdAddress[19] , GND_net);
    input sclk_c;
    output \port_status[19] ;
    output ws2813_out_c_19;
    input [23:0]\Q[19] ;
    output [8:0]\RdAddress[19] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1555;
    wire [31:0]n10927;
    
    wire sclk_c_enable_169, n54751, sclk_c_enable_170, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_173;
    wire [2:0]state_2__N_104;
    
    wire n14221, n53214, n53215;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53218, n53216, n53217, n53219, n54624, n54762, n54630, 
        n53373, n53374, n53375, n54851;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1373, n36543;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1365;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1404;
    wire [31:0]bit_counter_31__N_172;
    
    wire n54559;
    wire [31:0]n447;
    
    wire n54697;
    wire [31:0]n10751;
    
    wire n80, n14186, n54850, n42690;
    wire [8:0]n118;
    
    wire n53369, n53370, n53371, n53372, n54892, n54893, n54894, 
        n1, n1_adj_914, n71;
    wire [6:0]n15129;
    
    wire n10926, n52640, n37475, n42628, n4, n54629, n54567, n53206, 
        n53207, n54760;
    wire [31:0]n10853;
    
    wire n53208, n53209;
    wire [2:0]n6403;
    
    wire n36361, n53210, n53211, n53212, n53213, n53220, serial_N_437, 
        n36365, n6410;
    wire [31:0]bit_counter_31__N_204;
    
    wire n74, n48897, n48896, n48895, n48894, n48893, n48892, 
        n48891, n48890, n48889, n48888, n48887, n48886, n48885, 
        n48884, n48125, n48124, n48883, n48882, n48123, n48881, 
        n48880, n48879, n48878, n48877, n48876, n48875, n48874, 
        n48873, n48872, n48871, n48870, n48869, n48868, n48867, 
        n48866, n48122, n48121, n48120, n48119, n48118, n48117, 
        n48116, n48115, n48114, n47866, n47865, n48113, n48112, 
        n48111, n47864, n47863, n48110, n48108, n48107, n47862, 
        n48106, n47861, n47860, n48105, n47859, n47858, n47857, 
        n47856, n47855, n47854, n47853, n15, n14, n47852, n47851;
    
    FD1P3AX delay_counter_i0_i0 (.D(n10927[0]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54751), .SP(sclk_c_enable_169), .CK(sclk_c), 
            .Q(\port_status[19] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_170), .CK(sclk_c), 
            .Q(ws2813_out_c_19)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_173), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_173), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_173), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n14221), .Z(sclk_c_enable_173)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    L6MUX21 i38012 (.D0(n53214), .D1(n53215), .SD(bit_counter[2]), .Z(n53218));
    L6MUX21 i38013 (.D0(n53216), .D1(n53217), .SD(bit_counter[2]), .Z(n53219));
    LUT4 i1_2_lut_rep_621 (.A(state[1]), .B(n14221), .Z(n54624)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_621.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[1]), .B(n14221), .C(n54762), .D(n54630), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd080;
    L6MUX21 i38169 (.D0(n53373), .D1(n53374), .SD(bit_counter[2]), .Z(n53375));
    LUT4 i38471_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n14221), 
         .Z(n54851)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38471_4_lut_then_3_lut.init = 16'h1010;
    FD1P3IX pixel_i0 (.D(\Q[19] [0]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n54559), .B(n54762), .C(n447[8]), .D(n54697), 
         .Z(n10751[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_752 (.A(n54559), .B(n54762), .C(n447[12]), 
         .D(n54697), .Z(n10751[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_752.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_753 (.A(n54559), .B(n54762), .C(n447[9]), 
         .D(n54697), .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_753.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_754 (.A(n54559), .B(n54762), .C(n447[7]), 
         .D(n54697), .Z(n10751[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_754.init = 16'hf888;
    LUT4 i38471_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n14186), 
         .Z(n54850)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38471_4_lut_else_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n42690), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_755 (.A(state[2]), .B(n42690), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_755.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_756 (.A(state[2]), .B(n42690), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_756.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_757 (.A(state[2]), .B(n42690), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_757.init = 16'h1010;
    FD1P3AX delay_counter_i0_i1 (.D(n10927[1]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n10927[3]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_758 (.A(state[2]), .B(n42690), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_758.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_759 (.A(state[2]), .B(n42690), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_759.init = 16'h1010;
    FD1P3AX delay_counter_i0_i7 (.D(n10927[7]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n10927[8]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n10927[9]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_760 (.A(state[2]), .B(n42690), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_760.init = 16'h1010;
    FD1P3AX delay_counter_i0_i12 (.D(n10927[12]), .SP(sclk_c_enable_1555), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_761 (.A(state[2]), .B(n42690), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_761.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_762 (.A(state[2]), .B(n42690), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_762.init = 16'h1010;
    PFUMX i38167 (.BLUT(n53369), .ALUT(n53370), .C0(bit_counter[1]), .Z(n53373));
    PFUMX i38168 (.BLUT(n53371), .ALUT(n53372), .C0(bit_counter[1]), .Z(n53374));
    FD1P3IX pixel_i23 (.D(\Q[19] [23]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[19] [22]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[19] [21]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[19] [20]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[19] [19]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[19] [18]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[19] [17]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[19] [16]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[19] [15]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[19] [14]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[19] [13]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[19] [12]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[19] [11]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[19] [10]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[19] [9]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[19] [8]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[19] [7]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[19] [6]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[19] [5]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[19] [4]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[19] [3]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[19] [2]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[19] [1]), .SP(sclk_c_enable_1373), .CD(n36543), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1365), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1373), 
            .CD(n36543), .CK(sclk_c), .Q(\RdAddress[19] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    PFUMX i38903 (.BLUT(n54892), .ALUT(n54893), .C0(state[1]), .Z(n54894));
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1404), .CD(n36543), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_914), .SP(sclk_c_enable_1404), .CD(n36543), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1404), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 mux_2961_i2_4_lut (.A(n71), .B(n15129[0]), .C(n10926), .D(n52640), 
         .Z(n10927[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2961_i4_4_lut (.A(n37475), .B(n42628), .C(n10926), .D(n4), 
         .Z(n10927[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_3_lut_4_lut_4_lut_adj_763 (.A(n54762), .B(state[1]), .C(n54630), 
         .D(n54629), .Z(n52640)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_763.init = 16'hce02;
    LUT4 i1_4_lut (.A(n42690), .B(n54567), .C(n447[3]), .D(n54697), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    PFUMX i38008 (.BLUT(n53206), .ALUT(n53207), .C0(bit_counter[1]), .Z(n53214));
    LUT4 mux_2961_i8_4_lut (.A(n10751[7]), .B(n42628), .C(n10926), .D(n54567), 
         .Z(n10927[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i8_4_lut.init = 16'h303a;
    LUT4 mux_2951_i5_4_lut_4_lut (.A(state[0]), .B(n54760), .C(n447[4]), 
         .D(n54567), .Z(n10853[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2951_i5_4_lut_4_lut.init = 16'haad0;
    PFUMX i38009 (.BLUT(n53208), .ALUT(n53209), .C0(bit_counter[1]), .Z(n53215));
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n54760), .C(n14186), .D(n42690), 
         .Z(n6403[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfddd;
    LUT4 i24149_2_lut_4_lut (.A(n54629), .B(state[0]), .C(state[1]), .D(n10926), 
         .Z(n36361)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i24149_2_lut_4_lut.init = 16'hfd00;
    LUT4 mux_2961_i9_4_lut (.A(n10751[8]), .B(n42628), .C(n10926), .D(n54567), 
         .Z(n10927[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i9_4_lut.init = 16'h303a;
    LUT4 mux_2961_i10_4_lut (.A(n80), .B(n42628), .C(n10926), .D(n54567), 
         .Z(n10927[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i10_4_lut.init = 16'h303a;
    LUT4 mux_2961_i13_4_lut (.A(n10751[12]), .B(n42628), .C(n10926), .D(n54567), 
         .Z(n10927[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i13_4_lut.init = 16'h303a;
    PFUMX i38010 (.BLUT(n53210), .ALUT(n53211), .C0(bit_counter[1]), .Z(n53216));
    PFUMX i38011 (.BLUT(n53212), .ALUT(n53213), .C0(bit_counter[1]), .Z(n53217));
    LUT4 i38007_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38007_3_lut.init = 16'hcaca;
    LUT4 i38006_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38006_3_lut.init = 16'hcaca;
    LUT4 i38005_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38005_3_lut.init = 16'hcaca;
    LUT4 i38004_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38004_3_lut.init = 16'hcaca;
    LUT4 i38003_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38003_3_lut.init = 16'hcaca;
    LUT4 i38002_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38002_3_lut.init = 16'hcaca;
    LUT4 i38001_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38001_3_lut.init = 16'hcaca;
    LUT4 i38000_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38000_3_lut.init = 16'hcaca;
    LUT4 mux_2951_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14221), .Z(n54893)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2951_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2951_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14186), .Z(n54892)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2951_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53220), .B(n53375), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1555), 
            .CD(n36365), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1555), .CD(n36365), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1555), .CD(n36365), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n10853[4]), .SP(sclk_c_enable_1555), 
            .CD(n36361), .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54894), .SP(sclk_c_enable_1555), .CD(n36361), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=344, LSE_RLINE=344 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    L6MUX21 i38014 (.D0(n53218), .D1(n53219), .SD(bit_counter[3]), .Z(n53220));
    LUT4 i29446_4_lut (.A(n6403[0]), .B(n6410), .C(state[0]), .D(n54624), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29446_4_lut.init = 16'h0322;
    LUT4 i38166_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38166_3_lut.init = 16'hcaca;
    LUT4 i38165_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38165_3_lut.init = 16'hcaca;
    LUT4 i38164_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38164_3_lut.init = 16'hcaca;
    LUT4 i38163_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38163_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_764 (.A(state[2]), .B(state[0]), .C(state[1]), .D(n14221), 
         .Z(n6410)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_adj_764.init = 16'ha8a0;
    PFUMX i38875 (.BLUT(n54850), .ALUT(n54851), .C0(state[1]), .Z(state_2__N_104[1]));
    LUT4 i25266_1_lut_rep_748 (.A(state[2]), .Z(n54751)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25266_1_lut_rep_748.init = 16'h5555;
    LUT4 i29993_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i29993_3_lut_3_lut.init = 16'h5151;
    LUT4 i28794_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28794_2_lut.init = 16'hbbbb;
    LUT4 i38432_2_lut_rep_752 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1404)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38432_2_lut_rep_752.init = 16'h9999;
    LUT4 i28793_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_914)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28793_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_626 (.A(state[2]), .B(n14221), .Z(n54629)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_626.init = 16'h4444;
    LUT4 i1_2_lut_rep_757 (.A(state[1]), .B(state[2]), .Z(n54760)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_757.init = 16'heeee;
    LUT4 i1_2_lut_rep_694_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54697)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_694_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_765 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_765.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_766 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_766.init = 16'he0f0;
    LUT4 i24369_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36543)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i24369_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_767 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15129[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_767.init = 16'h7070;
    LUT4 i1_3_lut_rep_691_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1373)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_691_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n14221), 
         .Z(sclk_c_enable_170)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i30452_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42628)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i30452_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_759 (.A(state[0]), .B(state[2]), .Z(n54762)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_759.init = 16'h2222;
    LUT4 i1_2_lut_rep_564_3_lut (.A(state[2]), .B(n14221), .C(state[1]), 
         .Z(n54567)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_564_3_lut.init = 16'h4040;
    LUT4 i24173_4_lut (.A(sclk_c_enable_1555), .B(n54697), .C(n10926), 
         .D(n54567), .Z(n36365)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i24173_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_4_lut_adj_768 (.A(state[0]), .B(state[2]), .C(n14186), 
         .D(state[1]), .Z(n37475)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_768.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n14186), 
         .D(state[1]), .Z(sclk_c_enable_1365)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_769 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_769.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_770 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_770.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_771 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_771.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_772 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_772.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_773 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_773.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_774 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_774.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_775 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_775.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_776 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_776.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_777 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_777.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_778 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_778.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_779 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_779.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_780 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_780.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_781 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_781.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_782 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_782.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_783 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_783.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_784 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_784.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_785 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_785.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_786 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_786.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_787 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_787.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_788 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_788.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_789 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_789.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_790 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_790.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_791 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_791.init = 16'h2020;
    LUT4 i38572_3_lut_rep_565_4_lut (.A(state[2]), .B(n14221), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1555)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38572_3_lut_rep_565_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_adj_792 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_792.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_793 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_793.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_794 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_794.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_795 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_795.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_796 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_796.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_797 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_797.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_798 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_798.init = 16'h2020;
    LUT4 i1_2_lut_rep_627 (.A(n42690), .B(n14186), .Z(n54630)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_627.init = 16'h8888;
    LUT4 i1_2_lut_rep_556_3_lut (.A(n42690), .B(n14186), .C(state[1]), 
         .Z(n54559)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_556_3_lut.init = 16'h0808;
    CCU2D add_33932_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48897), 
          .S0(n14221));
    defparam add_33932_cout.INIT0 = 16'h0000;
    defparam add_33932_cout.INIT1 = 16'h0000;
    defparam add_33932_cout.INJECT1_0 = "NO";
    defparam add_33932_cout.INJECT1_1 = "NO";
    CCU2D add_33932_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48896), .COUT(n48897));
    defparam add_33932_31.INIT0 = 16'hf555;
    defparam add_33932_31.INIT1 = 16'h5555;
    defparam add_33932_31.INJECT1_0 = "NO";
    defparam add_33932_31.INJECT1_1 = "NO";
    CCU2D add_33932_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48895), .COUT(n48896));
    defparam add_33932_29.INIT0 = 16'hf555;
    defparam add_33932_29.INIT1 = 16'hf555;
    defparam add_33932_29.INJECT1_0 = "NO";
    defparam add_33932_29.INJECT1_1 = "NO";
    CCU2D add_33932_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48894), .COUT(n48895));
    defparam add_33932_27.INIT0 = 16'hf555;
    defparam add_33932_27.INIT1 = 16'hf555;
    defparam add_33932_27.INJECT1_0 = "NO";
    defparam add_33932_27.INJECT1_1 = "NO";
    CCU2D add_33932_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48893), .COUT(n48894));
    defparam add_33932_25.INIT0 = 16'hf555;
    defparam add_33932_25.INIT1 = 16'hf555;
    defparam add_33932_25.INJECT1_0 = "NO";
    defparam add_33932_25.INJECT1_1 = "NO";
    CCU2D add_33932_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48892), .COUT(n48893));
    defparam add_33932_23.INIT0 = 16'hf555;
    defparam add_33932_23.INIT1 = 16'hf555;
    defparam add_33932_23.INJECT1_0 = "NO";
    defparam add_33932_23.INJECT1_1 = "NO";
    CCU2D add_33932_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48891), .COUT(n48892));
    defparam add_33932_21.INIT0 = 16'hf555;
    defparam add_33932_21.INIT1 = 16'hf555;
    defparam add_33932_21.INJECT1_0 = "NO";
    defparam add_33932_21.INJECT1_1 = "NO";
    CCU2D add_33932_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48890), .COUT(n48891));
    defparam add_33932_19.INIT0 = 16'hf555;
    defparam add_33932_19.INIT1 = 16'hf555;
    defparam add_33932_19.INJECT1_0 = "NO";
    defparam add_33932_19.INJECT1_1 = "NO";
    CCU2D add_33932_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48889), .COUT(n48890));
    defparam add_33932_17.INIT0 = 16'hf555;
    defparam add_33932_17.INIT1 = 16'hf555;
    defparam add_33932_17.INJECT1_0 = "NO";
    defparam add_33932_17.INJECT1_1 = "NO";
    CCU2D add_33932_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48888), .COUT(n48889));
    defparam add_33932_15.INIT0 = 16'hf555;
    defparam add_33932_15.INIT1 = 16'hf555;
    defparam add_33932_15.INJECT1_0 = "NO";
    defparam add_33932_15.INJECT1_1 = "NO";
    CCU2D add_33932_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48887), .COUT(n48888));
    defparam add_33932_13.INIT0 = 16'hf555;
    defparam add_33932_13.INIT1 = 16'hf555;
    defparam add_33932_13.INJECT1_0 = "NO";
    defparam add_33932_13.INJECT1_1 = "NO";
    CCU2D add_33932_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48886), .COUT(n48887));
    defparam add_33932_11.INIT0 = 16'hf555;
    defparam add_33932_11.INIT1 = 16'hf555;
    defparam add_33932_11.INJECT1_0 = "NO";
    defparam add_33932_11.INJECT1_1 = "NO";
    CCU2D add_33932_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48885), .COUT(n48886));
    defparam add_33932_9.INIT0 = 16'hf555;
    defparam add_33932_9.INIT1 = 16'hf555;
    defparam add_33932_9.INJECT1_0 = "NO";
    defparam add_33932_9.INJECT1_1 = "NO";
    CCU2D add_33932_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48884), .COUT(n48885));
    defparam add_33932_7.INIT0 = 16'hf555;
    defparam add_33932_7.INIT1 = 16'hf555;
    defparam add_33932_7.INJECT1_0 = "NO";
    defparam add_33932_7.INJECT1_1 = "NO";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48125), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48124), .COUT(n48125), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_33932_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48883), .COUT(n48884));
    defparam add_33932_5.INIT0 = 16'hf555;
    defparam add_33932_5.INIT1 = 16'hf555;
    defparam add_33932_5.INJECT1_0 = "NO";
    defparam add_33932_5.INJECT1_1 = "NO";
    CCU2D add_33932_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48882), .COUT(n48883));
    defparam add_33932_3.INIT0 = 16'hf555;
    defparam add_33932_3.INIT1 = 16'hf555;
    defparam add_33932_3.INJECT1_0 = "NO";
    defparam add_33932_3.INJECT1_1 = "NO";
    CCU2D add_33932_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48882));
    defparam add_33932_1.INIT0 = 16'hF000;
    defparam add_33932_1.INIT1 = 16'ha666;
    defparam add_33932_1.INJECT1_0 = "NO";
    defparam add_33932_1.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48123), .COUT(n48124), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_33933_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48881), 
          .S0(n14186));
    defparam add_33933_cout.INIT0 = 16'h0000;
    defparam add_33933_cout.INIT1 = 16'h0000;
    defparam add_33933_cout.INJECT1_0 = "NO";
    defparam add_33933_cout.INJECT1_1 = "NO";
    CCU2D add_33933_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48880), .COUT(n48881));
    defparam add_33933_31.INIT0 = 16'hf555;
    defparam add_33933_31.INIT1 = 16'h5555;
    defparam add_33933_31.INJECT1_0 = "NO";
    defparam add_33933_31.INJECT1_1 = "NO";
    CCU2D add_33933_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48879), .COUT(n48880));
    defparam add_33933_29.INIT0 = 16'hf555;
    defparam add_33933_29.INIT1 = 16'hf555;
    defparam add_33933_29.INJECT1_0 = "NO";
    defparam add_33933_29.INJECT1_1 = "NO";
    CCU2D add_33933_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48878), .COUT(n48879));
    defparam add_33933_27.INIT0 = 16'hf555;
    defparam add_33933_27.INIT1 = 16'hf555;
    defparam add_33933_27.INJECT1_0 = "NO";
    defparam add_33933_27.INJECT1_1 = "NO";
    CCU2D add_33933_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48877), .COUT(n48878));
    defparam add_33933_25.INIT0 = 16'hf555;
    defparam add_33933_25.INIT1 = 16'hf555;
    defparam add_33933_25.INJECT1_0 = "NO";
    defparam add_33933_25.INJECT1_1 = "NO";
    CCU2D add_33933_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48876), .COUT(n48877));
    defparam add_33933_23.INIT0 = 16'hf555;
    defparam add_33933_23.INIT1 = 16'hf555;
    defparam add_33933_23.INJECT1_0 = "NO";
    defparam add_33933_23.INJECT1_1 = "NO";
    CCU2D add_33933_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48875), .COUT(n48876));
    defparam add_33933_21.INIT0 = 16'hf555;
    defparam add_33933_21.INIT1 = 16'hf555;
    defparam add_33933_21.INJECT1_0 = "NO";
    defparam add_33933_21.INJECT1_1 = "NO";
    CCU2D add_33933_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48874), .COUT(n48875));
    defparam add_33933_19.INIT0 = 16'hf555;
    defparam add_33933_19.INIT1 = 16'hf555;
    defparam add_33933_19.INJECT1_0 = "NO";
    defparam add_33933_19.INJECT1_1 = "NO";
    CCU2D add_33933_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48873), .COUT(n48874));
    defparam add_33933_17.INIT0 = 16'hf555;
    defparam add_33933_17.INIT1 = 16'hf555;
    defparam add_33933_17.INJECT1_0 = "NO";
    defparam add_33933_17.INJECT1_1 = "NO";
    CCU2D add_33933_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48872), .COUT(n48873));
    defparam add_33933_15.INIT0 = 16'hf555;
    defparam add_33933_15.INIT1 = 16'hf555;
    defparam add_33933_15.INJECT1_0 = "NO";
    defparam add_33933_15.INJECT1_1 = "NO";
    CCU2D add_33933_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48871), .COUT(n48872));
    defparam add_33933_13.INIT0 = 16'hf555;
    defparam add_33933_13.INIT1 = 16'hf555;
    defparam add_33933_13.INJECT1_0 = "NO";
    defparam add_33933_13.INJECT1_1 = "NO";
    CCU2D add_33933_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48870), .COUT(n48871));
    defparam add_33933_11.INIT0 = 16'hf555;
    defparam add_33933_11.INIT1 = 16'hf555;
    defparam add_33933_11.INJECT1_0 = "NO";
    defparam add_33933_11.INJECT1_1 = "NO";
    CCU2D add_33933_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48869), .COUT(n48870));
    defparam add_33933_9.INIT0 = 16'hf555;
    defparam add_33933_9.INIT1 = 16'hf555;
    defparam add_33933_9.INJECT1_0 = "NO";
    defparam add_33933_9.INJECT1_1 = "NO";
    CCU2D add_33933_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48868), .COUT(n48869));
    defparam add_33933_7.INIT0 = 16'hf555;
    defparam add_33933_7.INIT1 = 16'hf555;
    defparam add_33933_7.INJECT1_0 = "NO";
    defparam add_33933_7.INJECT1_1 = "NO";
    CCU2D add_33933_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48867), .COUT(n48868));
    defparam add_33933_5.INIT0 = 16'hf555;
    defparam add_33933_5.INIT1 = 16'hf555;
    defparam add_33933_5.INJECT1_0 = "NO";
    defparam add_33933_5.INJECT1_1 = "NO";
    CCU2D add_33933_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48866), .COUT(n48867));
    defparam add_33933_3.INIT0 = 16'hf555;
    defparam add_33933_3.INIT1 = 16'hf555;
    defparam add_33933_3.INJECT1_0 = "NO";
    defparam add_33933_3.INJECT1_1 = "NO";
    CCU2D add_33933_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48866));
    defparam add_33933_1.INIT0 = 16'hF000;
    defparam add_33933_1.INIT1 = 16'ha666;
    defparam add_33933_1.INJECT1_0 = "NO";
    defparam add_33933_1.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48122), .COUT(n48123), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48121), .COUT(n48122), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48120), .COUT(n48121), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48119), .COUT(n48120), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48118), .COUT(n48119), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48117), .COUT(n48118), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48116), .COUT(n48117), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48115), .COUT(n48116), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48114), .COUT(n48115), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_3140_33 (.A0(bit_counter[31]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47866), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_33.INIT0 = 16'h5999;
    defparam add_3140_33.INIT1 = 16'h0000;
    defparam add_3140_33.INJECT1_0 = "NO";
    defparam add_3140_33.INJECT1_1 = "NO";
    LUT4 mux_2961_i1_4_lut (.A(n74), .B(n15129[0]), .C(n10926), .D(n52640), 
         .Z(n10927[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2961_i1_4_lut.init = 16'hcfca;
    CCU2D add_3140_31 (.A0(bit_counter[29]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47865), .COUT(n47866), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_31.INIT0 = 16'h5999;
    defparam add_3140_31.INIT1 = 16'h5999;
    defparam add_3140_31.INJECT1_0 = "NO";
    defparam add_3140_31.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48113), .COUT(n48114), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48112), .COUT(n48113), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48111), .COUT(n48112), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_3140_29 (.A0(bit_counter[27]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47864), .COUT(n47865), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_29.INIT0 = 16'h5999;
    defparam add_3140_29.INIT1 = 16'h5999;
    defparam add_3140_29.INJECT1_0 = "NO";
    defparam add_3140_29.INJECT1_1 = "NO";
    CCU2D add_3140_27 (.A0(bit_counter[25]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47863), .COUT(n47864), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_27.INIT0 = 16'h5999;
    defparam add_3140_27.INIT1 = 16'h5999;
    defparam add_3140_27.INJECT1_0 = "NO";
    defparam add_3140_27.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48110), .COUT(n48111), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48110), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48108), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48107), .COUT(n48108), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_3140_25 (.A0(bit_counter[23]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47862), .COUT(n47863), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_25.INIT0 = 16'h5999;
    defparam add_3140_25.INIT1 = 16'h5999;
    defparam add_3140_25.INJECT1_0 = "NO";
    defparam add_3140_25.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48106), .COUT(n48107), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_3140_23 (.A0(bit_counter[21]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47861), .COUT(n47862), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_23.INIT0 = 16'h5999;
    defparam add_3140_23.INIT1 = 16'h5999;
    defparam add_3140_23.INJECT1_0 = "NO";
    defparam add_3140_23.INJECT1_1 = "NO";
    CCU2D add_3140_21 (.A0(bit_counter[19]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47860), .COUT(n47861), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_21.INIT0 = 16'h5999;
    defparam add_3140_21.INIT1 = 16'h5999;
    defparam add_3140_21.INJECT1_0 = "NO";
    defparam add_3140_21.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48105), .COUT(n48106), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48105), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3140_19 (.A0(bit_counter[17]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47859), .COUT(n47860), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_19.INIT0 = 16'h5999;
    defparam add_3140_19.INIT1 = 16'h5999;
    defparam add_3140_19.INJECT1_0 = "NO";
    defparam add_3140_19.INJECT1_1 = "NO";
    CCU2D add_3140_17 (.A0(bit_counter[15]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47858), .COUT(n47859), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_17.INIT0 = 16'h5999;
    defparam add_3140_17.INIT1 = 16'h5999;
    defparam add_3140_17.INJECT1_0 = "NO";
    defparam add_3140_17.INJECT1_1 = "NO";
    CCU2D add_3140_15 (.A0(bit_counter[13]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47857), .COUT(n47858), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_15.INIT0 = 16'h5999;
    defparam add_3140_15.INIT1 = 16'h5999;
    defparam add_3140_15.INJECT1_0 = "NO";
    defparam add_3140_15.INJECT1_1 = "NO";
    CCU2D add_3140_13 (.A0(bit_counter[11]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47856), .COUT(n47857), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_13.INIT0 = 16'h5999;
    defparam add_3140_13.INIT1 = 16'h5999;
    defparam add_3140_13.INJECT1_0 = "NO";
    defparam add_3140_13.INJECT1_1 = "NO";
    CCU2D add_3140_11 (.A0(bit_counter[9]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47855), .COUT(n47856), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_11.INIT0 = 16'h5999;
    defparam add_3140_11.INIT1 = 16'h5999;
    defparam add_3140_11.INJECT1_0 = "NO";
    defparam add_3140_11.INJECT1_1 = "NO";
    CCU2D add_3140_9 (.A0(bit_counter[7]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47854), .COUT(n47855), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_9.INIT0 = 16'h5999;
    defparam add_3140_9.INIT1 = 16'h5999;
    defparam add_3140_9.INJECT1_0 = "NO";
    defparam add_3140_9.INJECT1_1 = "NO";
    CCU2D add_3140_7 (.A0(bit_counter[5]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47853), .COUT(n47854), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_7.INIT0 = 16'h5999;
    defparam add_3140_7.INIT1 = 16'h5999;
    defparam add_3140_7.INJECT1_0 = "NO";
    defparam add_3140_7.INJECT1_1 = "NO";
    LUT4 i2973_3_lut (.A(state[2]), .B(state[1]), .C(n14221), .Z(n10926)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2973_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42690)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    CCU2D add_3140_5 (.A0(bit_counter[3]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47852), .COUT(n47853), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_5.INIT0 = 16'h5999;
    defparam add_3140_5.INIT1 = 16'h5999;
    defparam add_3140_5.INJECT1_0 = "NO";
    defparam add_3140_5.INJECT1_1 = "NO";
    CCU2D add_3140_3 (.A0(bit_counter[1]), .B0(n14186), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n14186), .C1(GND_net), 
          .D1(GND_net), .CIN(n47851), .COUT(n47852), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_3.INIT0 = 16'h5999;
    defparam add_3140_3.INIT1 = 16'h5999;
    defparam add_3140_3.INJECT1_0 = "NO";
    defparam add_3140_3.INJECT1_1 = "NO";
    CCU2D add_3140_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n14186), .C1(GND_net), .D1(GND_net), 
          .COUT(n47851), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3140_1.INIT0 = 16'hF000;
    defparam add_3140_1.INIT1 = 16'h5999;
    defparam add_3140_1.INJECT1_0 = "NO";
    defparam add_3140_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \spi_slave(8,'0','0','0') 
//

module \spi_slave(8,'0','0','0')  (rx_data_cnt, SCLK_SLAVE_c, rx_data_cnt_5__N_63, 
            n50005, sclk_c, RX_RDY, DATA_OUT, MOSI_SLAVE_c, CSn, 
            CSn_SLAVE_c, SCLK_SLAVE_c_enable_5);
    output [5:0]rx_data_cnt;
    input SCLK_SLAVE_c;
    output rx_data_cnt_5__N_63;
    input n50005;
    input sclk_c;
    output RX_RDY;
    output [7:0]DATA_OUT;
    input MOSI_SLAVE_c;
    input CSn;
    input CSn_SLAVE_c;
    input SCLK_SLAVE_c_enable_5;
    
    wire SCLK_SLAVE_c /* synthesis is_clock=1, SET_AS_NETWORK=SCLK_SLAVE_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(16[9:19])
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire rx_done, rx_done_flip1, rx_done_flip2, rx_done_flip3, n34110, 
        DATA_OUT_7__N_52;
    wire [7:0]rx_shift_data;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(76[13:26])
    
    wire CSn_SLAVE_N_56;
    wire [5:0]rx_data_cnt_c;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(91[25:36])
    
    wire n54785;
    wire [5:0]n90;
    
    wire n54708, n52913;
    
    FD1S3IX rx_data_cnt__i0 (.D(n50005), .CK(SCLK_SLAVE_c), .CD(rx_data_cnt_5__N_63), 
            .Q(rx_data_cnt[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i0.GSR = "ENABLED";
    FD1S3AX rx_done_145 (.D(rx_data_cnt_5__N_63), .CK(SCLK_SLAVE_c), .Q(rx_done)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(164[13] 172[20])
    defparam rx_done_145.GSR = "ENABLED";
    FD1S3AX rx_done_flip1_146 (.D(rx_done), .CK(sclk_c), .Q(rx_done_flip1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(301[6] 309[13])
    defparam rx_done_flip1_146.GSR = "ENABLED";
    FD1S3AX rx_done_flip2_147 (.D(rx_done_flip1), .CK(sclk_c), .Q(rx_done_flip2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(301[6] 309[13])
    defparam rx_done_flip2_147.GSR = "ENABLED";
    FD1S3AX rx_done_flip3_148 (.D(rx_done_flip2), .CK(sclk_c), .Q(rx_done_flip3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(301[6] 309[13])
    defparam rx_done_flip3_148.GSR = "ENABLED";
    FD1S3AX reg_rrdy_149 (.D(n34110), .CK(sclk_c), .Q(RX_RDY)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(314[6] 322[13])
    defparam reg_rrdy_149.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i0 (.D(rx_shift_data[0]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i0.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i0 (.D(MOSI_SLAVE_c), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i0.GSR = "ENABLED";
    LUT4 i21898_4_lut (.A(CSn), .B(rx_done_flip2), .C(RX_RDY), .D(rx_done_flip3), 
         .Z(n34110)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(314[6] 322[13])
    defparam i21898_4_lut.init = 16'ha0ec;
    LUT4 rx_done_flip1_I_0_2_lut (.A(rx_done_flip1), .B(rx_done_flip2), 
         .Z(DATA_OUT_7__N_52)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(117[12:51])
    defparam rx_done_flip1_I_0_2_lut.init = 16'h2222;
    LUT4 i3952_2_lut_rep_782 (.A(rx_data_cnt_c[1]), .B(rx_data_cnt[0]), 
         .Z(n54785)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3952_2_lut_rep_782.init = 16'h8888;
    LUT4 i3957_2_lut_3_lut (.A(rx_data_cnt_c[1]), .B(rx_data_cnt[0]), .C(rx_data_cnt_c[2]), 
         .Z(n90[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3957_2_lut_3_lut.init = 16'h7878;
    LUT4 i3959_2_lut_rep_705_3_lut (.A(rx_data_cnt_c[1]), .B(rx_data_cnt[0]), 
         .C(rx_data_cnt_c[2]), .Z(n54708)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3959_2_lut_rep_705_3_lut.init = 16'h8080;
    LUT4 i3964_2_lut_3_lut_4_lut (.A(rx_data_cnt_c[1]), .B(rx_data_cnt[0]), 
         .C(rx_data_cnt_c[3]), .D(rx_data_cnt_c[2]), .Z(n90[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3964_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 CSn_SLAVE_I_0_1_lut (.A(CSn_SLAVE_c), .Z(CSn_SLAVE_N_56)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(342[20:33])
    defparam CSn_SLAVE_I_0_1_lut.init = 16'h5555;
    FD1P3IX rx_data_cnt__i1 (.D(n90[1]), .SP(SCLK_SLAVE_c_enable_5), .CD(rx_data_cnt_5__N_63), 
            .CK(SCLK_SLAVE_c), .Q(rx_data_cnt_c[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i1.GSR = "ENABLED";
    FD1P3IX rx_data_cnt__i2 (.D(n90[2]), .SP(SCLK_SLAVE_c_enable_5), .CD(rx_data_cnt_5__N_63), 
            .CK(SCLK_SLAVE_c), .Q(rx_data_cnt_c[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i2.GSR = "ENABLED";
    FD1P3IX rx_data_cnt__i3 (.D(n90[3]), .SP(SCLK_SLAVE_c_enable_5), .CD(rx_data_cnt_5__N_63), 
            .CK(SCLK_SLAVE_c), .Q(rx_data_cnt_c[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i3.GSR = "ENABLED";
    FD1P3IX rx_data_cnt__i4 (.D(n90[4]), .SP(SCLK_SLAVE_c_enable_5), .CD(rx_data_cnt_5__N_63), 
            .CK(SCLK_SLAVE_c), .Q(rx_data_cnt_c[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i4.GSR = "ENABLED";
    FD1P3IX rx_data_cnt__i5 (.D(n90[5]), .SP(SCLK_SLAVE_c_enable_5), .CD(rx_data_cnt_5__N_63), 
            .CK(SCLK_SLAVE_c), .Q(rx_data_cnt_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(152[13] 160[20])
    defparam rx_data_cnt__i5.GSR = "ENABLED";
    LUT4 i38468_4_lut (.A(rx_data_cnt_c[3]), .B(rx_data_cnt_c[4]), .C(rx_data_cnt_c[5]), 
         .D(n52913), .Z(rx_data_cnt_5__N_63)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(155[19:48])
    defparam i38468_4_lut.init = 16'h0100;
    LUT4 i3978_3_lut_4_lut (.A(rx_data_cnt_c[3]), .B(n54708), .C(rx_data_cnt_c[4]), 
         .D(rx_data_cnt_c[5]), .Z(n90[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3978_3_lut_4_lut.init = 16'h7f80;
    FD1P3AX reg_rxdata_i0_i1 (.D(rx_shift_data[1]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i1.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i2 (.D(rx_shift_data[2]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i2.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i3 (.D(rx_shift_data[3]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i3.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i4 (.D(rx_shift_data[4]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i4.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i5 (.D(rx_shift_data[5]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i5.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i6 (.D(rx_shift_data[6]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i6.GSR = "ENABLED";
    FD1P3AX reg_rxdata_i0_i7 (.D(rx_shift_data[7]), .SP(DATA_OUT_7__N_52), 
            .CK(sclk_c), .Q(DATA_OUT[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(114[6] 120[13])
    defparam reg_rxdata_i0_i7.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i1 (.D(rx_shift_data[0]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i1.GSR = "ENABLED";
    LUT4 i3971_2_lut_3_lut_4_lut (.A(rx_data_cnt_c[2]), .B(n54785), .C(rx_data_cnt_c[4]), 
         .D(rx_data_cnt_c[3]), .Z(n90[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3971_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1P3AX rx_shift_data_i0_i2 (.D(rx_shift_data[1]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i2.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i3 (.D(rx_shift_data[2]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i3.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i4 (.D(rx_shift_data[3]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i4.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i5 (.D(rx_shift_data[4]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i5.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i6 (.D(rx_shift_data[5]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i6.GSR = "ENABLED";
    FD1P3AX rx_shift_data_i0_i7 (.D(rx_shift_data[6]), .SP(CSn_SLAVE_N_56), 
            .CK(SCLK_SLAVE_c), .Q(rx_shift_data[7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=21, LSE_LLINE=123, LSE_RLINE=123 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/simple_spi.vhd(138[13] 148[20])
    defparam rx_shift_data_i0_i7.GSR = "ENABLED";
    LUT4 i3950_2_lut (.A(rx_data_cnt_c[1]), .B(rx_data_cnt[0]), .Z(n90[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam i3950_2_lut.init = 16'h6666;
    LUT4 i37707_3_lut (.A(rx_data_cnt_c[1]), .B(rx_data_cnt_c[2]), .C(rx_data_cnt[0]), 
         .Z(n52913)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i37707_3_lut.init = 16'h8080;
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U33 
//

module \WS2812(48000000,"111111111")_U33  (sclk_c, \port_status[15] , ws2813_out_c_15, 
            \Q[15] , \RdAddress[15] , GND_net);
    input sclk_c;
    output \port_status[15] ;
    output ws2813_out_c_15;
    input [23:0]\Q[15] ;
    output [8:0]\RdAddress[15] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1935;
    wire [31:0]n9859;
    
    wire sclk_c_enable_138, n54768, sclk_c_enable_139, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_143;
    wire [2:0]state_2__N_104;
    
    wire n13941, n7488, n53154, n53155;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53158, n53156, n53157, n53159, n54641, n54584, n42682, 
        n13906, n54642, n54574, n54705;
    wire [31:0]n447;
    
    wire n103, n54962, n54961, n54779;
    wire [31:0]n9683;
    
    wire n76, n54859, n54860, n54861, n53345, n53346, n53347;
    wire [31:0]bit_counter_31__N_204;
    wire [31:0]bit_counter_31__N_172;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1753, n36163;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1720;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1784;
    wire [8:0]n118;
    
    wire n54700, n53146, n53147, n53148, n53149, n53150, n53151, 
        n53152, n53153, n53344, n53343, n53342, n53341, n52661, 
        n9858, n35981, n53160, n49150, n49149, n49148, n49147, 
        n49146, n49145, n49144, n49143, n49142, n49141, n49140, 
        n49139, n49138, n49137, n49136, n49135, n47967, n47966, 
        n47965, n47964, n47963, n47962, n36134, n47961, n47960, 
        n47959, n47958, n47957, n47956, n47955, n47954, n49054, 
        n47953, n49053, n49052, n49051, n49050, n49049, n49048, 
        n49047, n1, n1_adj_913, n49046, n49045, n49044, n49043, 
        n49042, n49041, n49040, n49039, n47952, n35985, n54963, 
        n69;
    wire [6:0]n15097;
    
    wire n15, n14, serial_N_437, n68, n38015, n4, n48041, n48040, 
        n48039, n48038, n48037, n48036, n48035, n48034, n48033, 
        n48032, n48031, n48030, n48029, n48028, n48027, n48026, 
        n48024, n48023, n48022, n48021;
    
    FD1P3AX delay_counter_i0_i0 (.D(n9859[0]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54768), .SP(sclk_c_enable_138), .CK(sclk_c), 
            .Q(\port_status[15] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_139), .CK(sclk_c), 
            .Q(ws2813_out_c_15)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_143), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_143), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_143), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13941), .Z(n7488)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 i38464_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13941), .Z(sclk_c_enable_143)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38464_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    L6MUX21 i37952 (.D0(n53154), .D1(n53155), .SD(bit_counter[2]), .Z(n53158));
    L6MUX21 i37953 (.D0(n53156), .D1(n53157), .SD(bit_counter[2]), .Z(n53159));
    LUT4 i1_2_lut_rep_638 (.A(state[2]), .B(n13941), .Z(n54641)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_638.init = 16'h4444;
    LUT4 i1_2_lut_rep_581_3_lut (.A(state[2]), .B(n13941), .C(state[1]), 
         .Z(n54584)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_581_3_lut.init = 16'h4040;
    LUT4 i38580_3_lut_rep_583_4_lut (.A(state[2]), .B(n13941), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1935)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38580_3_lut_rep_583_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_rep_639 (.A(n42682), .B(n13906), .Z(n54642)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_639.init = 16'h8888;
    LUT4 i1_2_lut_rep_571_3_lut (.A(n42682), .B(n13906), .C(state[1]), 
         .Z(n54574)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_571_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42682), .B(n13906), .C(n54705), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2723_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13941), .Z(n54962)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2723_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2723_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13941), .Z(n54961)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2723_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 i1_3_lut_4_lut (.A(n54574), .B(n54779), .C(n447[7]), .D(n54705), 
         .Z(n9683[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_709 (.A(n54574), .B(n54779), .C(n447[8]), 
         .D(n54705), .Z(n9683[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_709.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_710 (.A(n54574), .B(n54779), .C(n447[9]), 
         .D(n54705), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_710.init = 16'hf888;
    PFUMX i38881 (.BLUT(n54859), .ALUT(n54860), .C0(state[1]), .Z(n54861));
    L6MUX21 i38141 (.D0(n53345), .D1(n53346), .SD(bit_counter[2]), .Z(n53347));
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    FD1P3IX pixel_i0 (.D(\Q[15] [0]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i1 (.D(n9859[1]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n9859[3]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n9859[7]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n9859[8]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n9859[9]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n9859[12]), .SP(sclk_c_enable_1935), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_711 (.A(state[2]), .B(n42682), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_711.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_712 (.A(state[2]), .B(n42682), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_712.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_713 (.A(state[2]), .B(n42682), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_713.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_714 (.A(state[2]), .B(n42682), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_714.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_715 (.A(state[2]), .B(n42682), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_715.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_716 (.A(state[2]), .B(n42682), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_716.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_717 (.A(state[2]), .B(n42682), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_717.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_718 (.A(state[2]), .B(n42682), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_718.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_719 (.A(state[2]), .B(n42682), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_719.init = 16'h1010;
    LUT4 mux_2224_i2_4_lut_4_lut (.A(n54700), .B(n54705), .C(n7488), .D(n13906), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2224_i2_4_lut_4_lut.init = 16'h5053;
    PFUMX i37948 (.BLUT(n53146), .ALUT(n53147), .C0(bit_counter[1]), .Z(n53154));
    LUT4 i1_2_lut_3_lut_adj_720 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_720.init = 16'h2020;
    PFUMX i37949 (.BLUT(n53148), .ALUT(n53149), .C0(bit_counter[1]), .Z(n53155));
    PFUMX i37950 (.BLUT(n53150), .ALUT(n53151), .C0(bit_counter[1]), .Z(n53156));
    PFUMX i37951 (.BLUT(n53152), .ALUT(n53153), .C0(bit_counter[1]), .Z(n53157));
    LUT4 i38138_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38138_3_lut.init = 16'hcaca;
    LUT4 i38137_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38137_3_lut.init = 16'hcaca;
    LUT4 i38136_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38136_3_lut.init = 16'hcaca;
    LUT4 i38135_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38135_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54642), .C(n13941), .D(n54779), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54779), .B(state[1]), .C(n54642), .D(n54641), 
         .Z(n52661)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 i23769_2_lut_4_lut (.A(n54641), .B(state[0]), .C(state[1]), .D(n9858), 
         .Z(n35981)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23769_2_lut_4_lut.init = 16'hfd00;
    LUT4 i1_2_lut_3_lut_adj_721 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_721.init = 16'h2020;
    LUT4 i37947_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37947_3_lut.init = 16'hcaca;
    LUT4 i37946_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37946_3_lut.init = 16'hcaca;
    LUT4 i37945_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37945_3_lut.init = 16'hcaca;
    LUT4 i37944_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37944_3_lut.init = 16'hcaca;
    LUT4 i37943_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37943_3_lut.init = 16'hcaca;
    LUT4 i37942_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37942_3_lut.init = 16'hcaca;
    LUT4 i37941_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37941_3_lut.init = 16'hcaca;
    LUT4 i37940_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37940_3_lut.init = 16'hcaca;
    L6MUX21 i37954 (.D0(n53158), .D1(n53159), .SD(bit_counter[3]), .Z(n53160));
    CCU2D add_33900_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49150), 
          .S0(n13941));
    defparam add_33900_cout.INIT0 = 16'h0000;
    defparam add_33900_cout.INIT1 = 16'h0000;
    defparam add_33900_cout.INJECT1_0 = "NO";
    defparam add_33900_cout.INJECT1_1 = "NO";
    CCU2D add_33900_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49149), .COUT(n49150));
    defparam add_33900_31.INIT0 = 16'hf555;
    defparam add_33900_31.INIT1 = 16'h5555;
    defparam add_33900_31.INJECT1_0 = "NO";
    defparam add_33900_31.INJECT1_1 = "NO";
    CCU2D add_33900_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49148), .COUT(n49149));
    defparam add_33900_29.INIT0 = 16'hf555;
    defparam add_33900_29.INIT1 = 16'hf555;
    defparam add_33900_29.INJECT1_0 = "NO";
    defparam add_33900_29.INJECT1_1 = "NO";
    CCU2D add_33900_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49147), .COUT(n49148));
    defparam add_33900_27.INIT0 = 16'hf555;
    defparam add_33900_27.INIT1 = 16'hf555;
    defparam add_33900_27.INJECT1_0 = "NO";
    defparam add_33900_27.INJECT1_1 = "NO";
    PFUMX i38139 (.BLUT(n53341), .ALUT(n53342), .C0(bit_counter[1]), .Z(n53345));
    CCU2D add_33900_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49146), .COUT(n49147));
    defparam add_33900_25.INIT0 = 16'hf555;
    defparam add_33900_25.INIT1 = 16'hf555;
    defparam add_33900_25.INJECT1_0 = "NO";
    defparam add_33900_25.INJECT1_1 = "NO";
    CCU2D add_33900_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49145), .COUT(n49146));
    defparam add_33900_23.INIT0 = 16'hf555;
    defparam add_33900_23.INIT1 = 16'hf555;
    defparam add_33900_23.INJECT1_0 = "NO";
    defparam add_33900_23.INJECT1_1 = "NO";
    CCU2D add_33900_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49144), .COUT(n49145));
    defparam add_33900_21.INIT0 = 16'hf555;
    defparam add_33900_21.INIT1 = 16'hf555;
    defparam add_33900_21.INJECT1_0 = "NO";
    defparam add_33900_21.INJECT1_1 = "NO";
    CCU2D add_33900_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49143), .COUT(n49144));
    defparam add_33900_19.INIT0 = 16'hf555;
    defparam add_33900_19.INIT1 = 16'hf555;
    defparam add_33900_19.INJECT1_0 = "NO";
    defparam add_33900_19.INJECT1_1 = "NO";
    CCU2D add_33900_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49142), .COUT(n49143));
    defparam add_33900_17.INIT0 = 16'hf555;
    defparam add_33900_17.INIT1 = 16'hf555;
    defparam add_33900_17.INJECT1_0 = "NO";
    defparam add_33900_17.INJECT1_1 = "NO";
    CCU2D add_33900_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49141), .COUT(n49142));
    defparam add_33900_15.INIT0 = 16'hf555;
    defparam add_33900_15.INIT1 = 16'hf555;
    defparam add_33900_15.INJECT1_0 = "NO";
    defparam add_33900_15.INJECT1_1 = "NO";
    CCU2D add_33900_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49140), .COUT(n49141));
    defparam add_33900_13.INIT0 = 16'hf555;
    defparam add_33900_13.INIT1 = 16'hf555;
    defparam add_33900_13.INJECT1_0 = "NO";
    defparam add_33900_13.INJECT1_1 = "NO";
    CCU2D add_33900_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49139), .COUT(n49140));
    defparam add_33900_11.INIT0 = 16'hf555;
    defparam add_33900_11.INIT1 = 16'hf555;
    defparam add_33900_11.INJECT1_0 = "NO";
    defparam add_33900_11.INJECT1_1 = "NO";
    CCU2D add_33900_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49138), .COUT(n49139));
    defparam add_33900_9.INIT0 = 16'hf555;
    defparam add_33900_9.INIT1 = 16'hf555;
    defparam add_33900_9.INJECT1_0 = "NO";
    defparam add_33900_9.INJECT1_1 = "NO";
    CCU2D add_33900_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49137), .COUT(n49138));
    defparam add_33900_7.INIT0 = 16'hf555;
    defparam add_33900_7.INIT1 = 16'hf555;
    defparam add_33900_7.INJECT1_0 = "NO";
    defparam add_33900_7.INJECT1_1 = "NO";
    CCU2D add_33900_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49136), .COUT(n49137));
    defparam add_33900_5.INIT0 = 16'hf555;
    defparam add_33900_5.INIT1 = 16'hf555;
    defparam add_33900_5.INJECT1_0 = "NO";
    defparam add_33900_5.INJECT1_1 = "NO";
    CCU2D add_33900_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49135), .COUT(n49136));
    defparam add_33900_3.INIT0 = 16'hf555;
    defparam add_33900_3.INIT1 = 16'hf555;
    defparam add_33900_3.INJECT1_0 = "NO";
    defparam add_33900_3.INJECT1_1 = "NO";
    PFUMX i38140 (.BLUT(n53343), .ALUT(n53344), .C0(bit_counter[1]), .Z(n53346));
    CCU2D add_33900_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n49135));
    defparam add_33900_1.INIT0 = 16'hF000;
    defparam add_33900_1.INIT1 = 16'ha666;
    defparam add_33900_1.INJECT1_0 = "NO";
    defparam add_33900_1.INJECT1_1 = "NO";
    CCU2D add_3132_33 (.A0(bit_counter[31]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47967), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_33.INIT0 = 16'h5999;
    defparam add_3132_33.INIT1 = 16'h0000;
    defparam add_3132_33.INJECT1_0 = "NO";
    defparam add_3132_33.INJECT1_1 = "NO";
    CCU2D add_3132_31 (.A0(bit_counter[29]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47966), .COUT(n47967), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_31.INIT0 = 16'h5999;
    defparam add_3132_31.INIT1 = 16'h5999;
    defparam add_3132_31.INJECT1_0 = "NO";
    defparam add_3132_31.INJECT1_1 = "NO";
    CCU2D add_3132_29 (.A0(bit_counter[27]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47965), .COUT(n47966), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_29.INIT0 = 16'h5999;
    defparam add_3132_29.INIT1 = 16'h5999;
    defparam add_3132_29.INJECT1_0 = "NO";
    defparam add_3132_29.INJECT1_1 = "NO";
    CCU2D add_3132_27 (.A0(bit_counter[25]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47964), .COUT(n47965), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_27.INIT0 = 16'h5999;
    defparam add_3132_27.INIT1 = 16'h5999;
    defparam add_3132_27.INJECT1_0 = "NO";
    defparam add_3132_27.INJECT1_1 = "NO";
    CCU2D add_3132_25 (.A0(bit_counter[23]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47963), .COUT(n47964), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_25.INIT0 = 16'h5999;
    defparam add_3132_25.INIT1 = 16'h5999;
    defparam add_3132_25.INJECT1_0 = "NO";
    defparam add_3132_25.INJECT1_1 = "NO";
    FD1P3IX pixel_i23 (.D(\Q[15] [23]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[15] [22]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    CCU2D add_3132_23 (.A0(bit_counter[21]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47962), .COUT(n47963), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_23.INIT0 = 16'h5999;
    defparam add_3132_23.INIT1 = 16'h5999;
    defparam add_3132_23.INJECT1_0 = "NO";
    defparam add_3132_23.INJECT1_1 = "NO";
    FD1P3IX pixel_i21 (.D(\Q[15] [21]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[15] [20]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[15] [19]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[15] [18]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[15] [17]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    LUT4 i38418_2_lut_rep_742 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1784)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38418_2_lut_rep_742.init = 16'h9999;
    FD1P3IX pixel_i16 (.D(\Q[15] [16]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[15] [15]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    LUT4 i23922_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36134)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23922_2_lut_2_lut.init = 16'h8888;
    FD1P3IX pixel_i14 (.D(\Q[15] [14]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[15] [13]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[15] [12]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[15] [11]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[15] [10]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[15] [9]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[15] [8]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[15] [7]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[15] [6]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[15] [5]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[15] [4]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[15] [3]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[15] [2]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[15] [1]), .SP(sclk_c_enable_1753), .CD(n36163), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    CCU2D add_3132_21 (.A0(bit_counter[19]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47961), .COUT(n47962), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_21.INIT0 = 16'h5999;
    defparam add_3132_21.INIT1 = 16'h5999;
    defparam add_3132_21.INJECT1_0 = "NO";
    defparam add_3132_21.INJECT1_1 = "NO";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1720), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    CCU2D add_3132_19 (.A0(bit_counter[17]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47960), .COUT(n47961), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_19.INIT0 = 16'h5999;
    defparam add_3132_19.INIT1 = 16'h5999;
    defparam add_3132_19.INJECT1_0 = "NO";
    defparam add_3132_19.INJECT1_1 = "NO";
    CCU2D add_3132_17 (.A0(bit_counter[15]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47959), .COUT(n47960), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_17.INIT0 = 16'h5999;
    defparam add_3132_17.INIT1 = 16'h5999;
    defparam add_3132_17.INJECT1_0 = "NO";
    defparam add_3132_17.INJECT1_1 = "NO";
    CCU2D add_3132_15 (.A0(bit_counter[13]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47958), .COUT(n47959), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_15.INIT0 = 16'h5999;
    defparam add_3132_15.INIT1 = 16'h5999;
    defparam add_3132_15.INJECT1_0 = "NO";
    defparam add_3132_15.INJECT1_1 = "NO";
    CCU2D add_3132_13 (.A0(bit_counter[11]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47957), .COUT(n47958), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_13.INIT0 = 16'h5999;
    defparam add_3132_13.INIT1 = 16'h5999;
    defparam add_3132_13.INJECT1_0 = "NO";
    defparam add_3132_13.INJECT1_1 = "NO";
    CCU2D add_3132_11 (.A0(bit_counter[9]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47956), .COUT(n47957), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_11.INIT0 = 16'h5999;
    defparam add_3132_11.INIT1 = 16'h5999;
    defparam add_3132_11.INJECT1_0 = "NO";
    defparam add_3132_11.INJECT1_1 = "NO";
    CCU2D add_3132_9 (.A0(bit_counter[7]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47955), .COUT(n47956), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_9.INIT0 = 16'h5999;
    defparam add_3132_9.INIT1 = 16'h5999;
    defparam add_3132_9.INJECT1_0 = "NO";
    defparam add_3132_9.INJECT1_1 = "NO";
    CCU2D add_3132_7 (.A0(bit_counter[5]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47954), .COUT(n47955), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_7.INIT0 = 16'h5999;
    defparam add_3132_7.INIT1 = 16'h5999;
    defparam add_3132_7.INJECT1_0 = "NO";
    defparam add_3132_7.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1753), 
            .CD(n36163), .CK(sclk_c), .Q(\RdAddress[15] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    CCU2D add_33901_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49054), 
          .S0(n13906));
    defparam add_33901_cout.INIT0 = 16'h0000;
    defparam add_33901_cout.INIT1 = 16'h0000;
    defparam add_33901_cout.INJECT1_0 = "NO";
    defparam add_33901_cout.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    CCU2D add_3132_5 (.A0(bit_counter[3]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47953), .COUT(n47954), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_5.INIT0 = 16'h5999;
    defparam add_3132_5.INIT1 = 16'h5999;
    defparam add_3132_5.INJECT1_0 = "NO";
    defparam add_3132_5.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    CCU2D add_33901_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49053), .COUT(n49054));
    defparam add_33901_31.INIT0 = 16'hf555;
    defparam add_33901_31.INIT1 = 16'h5555;
    defparam add_33901_31.INJECT1_0 = "NO";
    defparam add_33901_31.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    CCU2D add_33901_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49052), .COUT(n49053));
    defparam add_33901_29.INIT0 = 16'hf555;
    defparam add_33901_29.INIT1 = 16'hf555;
    defparam add_33901_29.INJECT1_0 = "NO";
    defparam add_33901_29.INJECT1_1 = "NO";
    CCU2D add_33901_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49051), .COUT(n49052));
    defparam add_33901_27.INIT0 = 16'hf555;
    defparam add_33901_27.INIT1 = 16'hf555;
    defparam add_33901_27.INJECT1_0 = "NO";
    defparam add_33901_27.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    CCU2D add_33901_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49050), .COUT(n49051));
    defparam add_33901_25.INIT0 = 16'hf555;
    defparam add_33901_25.INIT1 = 16'hf555;
    defparam add_33901_25.INJECT1_0 = "NO";
    defparam add_33901_25.INJECT1_1 = "NO";
    CCU2D add_33901_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49049), .COUT(n49050));
    defparam add_33901_23.INIT0 = 16'hf555;
    defparam add_33901_23.INIT1 = 16'hf555;
    defparam add_33901_23.INJECT1_0 = "NO";
    defparam add_33901_23.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    CCU2D add_33901_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49048), .COUT(n49049));
    defparam add_33901_21.INIT0 = 16'hf555;
    defparam add_33901_21.INIT1 = 16'hf555;
    defparam add_33901_21.INJECT1_0 = "NO";
    defparam add_33901_21.INJECT1_1 = "NO";
    CCU2D add_33901_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49047), .COUT(n49048));
    defparam add_33901_19.INIT0 = 16'hf555;
    defparam add_33901_19.INIT1 = 16'hf555;
    defparam add_33901_19.INJECT1_0 = "NO";
    defparam add_33901_19.INJECT1_1 = "NO";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1784), .CD(n36134), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_913), .SP(sclk_c_enable_1784), .CD(n36134), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    CCU2D add_33901_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49046), .COUT(n49047));
    defparam add_33901_17.INIT0 = 16'hf555;
    defparam add_33901_17.INIT1 = 16'hf555;
    defparam add_33901_17.INJECT1_0 = "NO";
    defparam add_33901_17.INJECT1_1 = "NO";
    CCU2D add_33901_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49045), .COUT(n49046));
    defparam add_33901_15.INIT0 = 16'hf555;
    defparam add_33901_15.INIT1 = 16'hf555;
    defparam add_33901_15.INJECT1_0 = "NO";
    defparam add_33901_15.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    CCU2D add_33901_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49044), .COUT(n49045));
    defparam add_33901_13.INIT0 = 16'hf555;
    defparam add_33901_13.INIT1 = 16'hf555;
    defparam add_33901_13.INJECT1_0 = "NO";
    defparam add_33901_13.INJECT1_1 = "NO";
    CCU2D add_33901_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49043), .COUT(n49044));
    defparam add_33901_11.INIT0 = 16'hf555;
    defparam add_33901_11.INIT1 = 16'hf555;
    defparam add_33901_11.INJECT1_0 = "NO";
    defparam add_33901_11.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1784), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    CCU2D add_33901_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49042), .COUT(n49043));
    defparam add_33901_9.INIT0 = 16'hf555;
    defparam add_33901_9.INIT1 = 16'hf555;
    defparam add_33901_9.INJECT1_0 = "NO";
    defparam add_33901_9.INJECT1_1 = "NO";
    CCU2D add_33901_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49041), .COUT(n49042));
    defparam add_33901_7.INIT0 = 16'hf555;
    defparam add_33901_7.INIT1 = 16'hf555;
    defparam add_33901_7.INJECT1_0 = "NO";
    defparam add_33901_7.INJECT1_1 = "NO";
    CCU2D add_33901_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49040), .COUT(n49041));
    defparam add_33901_5.INIT0 = 16'hf555;
    defparam add_33901_5.INIT1 = 16'hf555;
    defparam add_33901_5.INJECT1_0 = "NO";
    defparam add_33901_5.INJECT1_1 = "NO";
    CCU2D add_33901_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49039), .COUT(n49040));
    defparam add_33901_3.INIT0 = 16'hf555;
    defparam add_33901_3.INIT1 = 16'hf555;
    defparam add_33901_3.INJECT1_0 = "NO";
    defparam add_33901_3.INJECT1_1 = "NO";
    CCU2D add_33901_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n49039));
    defparam add_33901_1.INIT0 = 16'hF000;
    defparam add_33901_1.INIT1 = 16'ha666;
    defparam add_33901_1.INJECT1_0 = "NO";
    defparam add_33901_1.INJECT1_1 = "NO";
    CCU2D add_3132_3 (.A0(bit_counter[1]), .B0(n13906), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13906), .C1(GND_net), 
          .D1(GND_net), .CIN(n47952), .COUT(n47953), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_3.INIT0 = 16'h5999;
    defparam add_3132_3.INIT1 = 16'h5999;
    defparam add_3132_3.INJECT1_0 = "NO";
    defparam add_3132_3.INJECT1_1 = "NO";
    CCU2D add_3132_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13906), .C1(GND_net), .D1(GND_net), 
          .COUT(n47952), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3132_1.INIT0 = 16'hF000;
    defparam add_3132_1.INIT1 = 16'h5999;
    defparam add_3132_1.INJECT1_0 = "NO";
    defparam add_3132_1.INJECT1_1 = "NO";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1935), 
            .CD(n35985), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1935), .CD(n35985), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1935), .CD(n35985), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54963), .SP(sclk_c_enable_1935), .CD(n35981), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54861), .SP(sclk_c_enable_1935), .CD(n35981), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=300, LSE_RLINE=300 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_697_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54700)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_697_3_lut.init = 16'hf8f8;
    LUT4 mux_2733_i1_4_lut (.A(n69), .B(n15097[0]), .C(n9858), .D(n52661), 
         .Z(n9859[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i1_4_lut.init = 16'hcfca;
    LUT4 i2745_3_lut (.A(state[2]), .B(state[1]), .C(n13941), .Z(n9858)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2745_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42682)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 mux_2723_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13941), .Z(n54860)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2723_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2723_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13906), .Z(n54859)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2723_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53160), .B(n53347), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_3_lut_adj_722 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_722.init = 16'h2020;
    LUT4 mux_2224_i1_4_lut (.A(n54642), .B(n54700), .C(n7488), .D(n54705), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2224_i1_4_lut.init = 16'h3f3a;
    LUT4 i1_2_lut_3_lut_adj_723 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15097[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_723.init = 16'h7070;
    LUT4 i1_2_lut_rep_702_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54705)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_702_3_lut.init = 16'hefef;
    LUT4 i25813_1_lut_rep_765 (.A(state[2]), .Z(n54768)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25813_1_lut_rep_765.init = 16'h5555;
    LUT4 i28952_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28952_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n13941), 
         .Z(sclk_c_enable_139)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i28786_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28786_2_lut.init = 16'hbbbb;
    LUT4 i28785_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_913)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28785_2_lut.init = 16'hbbbb;
    LUT4 i1_3_lut_rep_684_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_1753)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_684_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_724 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_724.init = 16'he0f0;
    LUT4 i24014_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n36163)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i24014_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_776 (.A(state[0]), .B(state[2]), .Z(n54779)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_776.init = 16'h2222;
    LUT4 mux_2733_i2_4_lut (.A(n68), .B(n15097[0]), .C(n9858), .D(n52661), 
         .Z(n9859[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i2_4_lut.init = 16'hcfca;
    LUT4 i23793_4_lut (.A(sclk_c_enable_1935), .B(n54705), .C(n9858), 
         .D(n54584), .Z(n35985)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23793_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_4_lut_adj_725 (.A(state[0]), .B(state[2]), .C(n13906), 
         .D(state[1]), .Z(n38015)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_725.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_adj_726 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_726.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_727 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_727.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_728 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_728.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13906), 
         .D(state[1]), .Z(sclk_c_enable_1720)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_729 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_729.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_730 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_730.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_731 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_731.init = 16'h2020;
    LUT4 mux_2733_i4_4_lut (.A(n38015), .B(n54700), .C(n9858), .D(n4), 
         .Z(n9859[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_2_lut_3_lut_adj_732 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_732.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_733 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_733.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_734 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_734.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_735 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_735.init = 16'h2020;
    LUT4 mux_2733_i10_4_lut (.A(n76), .B(n54700), .C(n9858), .D(n54584), 
         .Z(n9859[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i10_4_lut.init = 16'h303a;
    LUT4 i1_2_lut_3_lut_adj_736 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_736.init = 16'h2020;
    LUT4 i1_4_lut (.A(n42682), .B(n54584), .C(n447[3]), .D(n54705), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2733_i13_4_lut (.A(n54584), .B(n54700), .C(n9858), .D(n103), 
         .Z(n9859[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i13_4_lut.init = 16'h3530;
    LUT4 i1_2_lut_3_lut_adj_737 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_737.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_738 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_738.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_739 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_739.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_740 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_740.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_741 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_741.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_742 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_742.init = 16'h2020;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48041), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    LUT4 mux_2733_i8_4_lut (.A(n9683[7]), .B(n54700), .C(n9858), .D(n54584), 
         .Z(n9859[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i8_4_lut.init = 16'h303a;
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48040), .COUT(n48041), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48039), .COUT(n48040), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48038), .COUT(n48039), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48037), .COUT(n48038), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48036), .COUT(n48037), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48035), .COUT(n48036), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48034), .COUT(n48035), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_743 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_743.init = 16'h2020;
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48033), .COUT(n48034), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_744 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_744.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_745 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_745.init = 16'h2020;
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48032), .COUT(n48033), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48031), .COUT(n48032), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    LUT4 mux_2733_i9_4_lut (.A(n9683[8]), .B(n54700), .C(n9858), .D(n54584), 
         .Z(n9859[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2733_i9_4_lut.init = 16'h303a;
    LUT4 i1_2_lut_3_lut_adj_746 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_746.init = 16'h2020;
    PFUMX i38949 (.BLUT(n54961), .ALUT(n54962), .C0(state[0]), .Z(n54963));
    LUT4 i1_2_lut_3_lut_adj_747 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_747.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_748 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_748.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_749 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_749.init = 16'h2020;
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48030), .COUT(n48031), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48029), .COUT(n48030), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_750 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_750.init = 16'h2020;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48028), .COUT(n48029), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_751 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_751.init = 16'h2020;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48027), .COUT(n48028), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48026), .COUT(n48027), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48026), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48024), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48023), .COUT(n48024), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48022), .COUT(n48023), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48021), .COUT(n48022), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48021), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U31 
//

module \WS2812(48000000,"111111111")_U31  (sclk_c, \port_status[17] , ws2813_out_c_17, 
            \Q[17] , \RdAddress[17] , GND_net);
    input sclk_c;
    output \port_status[17] ;
    output ws2813_out_c_17;
    input [23:0]\Q[17] ;
    output [8:0]\RdAddress[17] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1745;
    wire [31:0]n10393;
    
    wire sclk_c_enable_154, n54759, sclk_c_enable_155, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_158;
    wire [2:0]state_2__N_104;
    
    wire n14081, n6954, n14046, sclk_c_enable_1530, n53184, n53185;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53188, n53186, n53187, n53189;
    wire [31:0]n447;
    
    wire n54968, n54967, n54872, n54871, n53359, n53360, n53361, 
        n68;
    wire [6:0]n15113;
    
    wire n10392, n52664, n37745, n54696, n4, n42686, n54576, n54701;
    wire [31:0]n10217;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1563, n36353;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1594;
    wire [31:0]bit_counter_31__N_172;
    
    wire n76, n103;
    wire [8:0]n118;
    
    wire n54565, n54770, n53176, n53177, n53358, n53178, n53179, 
        n53357, n53356, n53180, n53181, n53355, n53182, n53183, 
        n54636, n54635, n36171, n53190, n1, n1_adj_912, n36175, 
        n54969, n54873, n47935;
    wire [31:0]bit_counter_31__N_204;
    
    wire n47934, n47933, n47932, n47931, n47930, n47929, n47928, 
        n47927, serial_N_437, n47926, n47925, n47924, n47923, n47922, 
        n47921, n47920, n69, n15, n14, n48083, n48082, n48081, 
        n48080, n48079, n48078, n48077, n48076, n48075, n48074, 
        n48073, n48072, n48071, n48070, n48069, n48068, n48721, 
        n48720, n48719, n48718, n48717, n48716, n48715, n48714, 
        n48713, n48712, n48066, n48065, n48711, n48710, n48709, 
        n48708, n48707, n48706, n48064, n48063, n48625, n48624, 
        n48623, n48622, n48621, n48620, n48619, n48618, n48617, 
        n48616, n48615, n48614, n48613, n48612, n48611, n48610;
    
    FD1P3AX delay_counter_i0_i0 (.D(n10393[0]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54759), .SP(sclk_c_enable_154), .CK(sclk_c), 
            .Q(\port_status[17] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_155), .CK(sclk_c), 
            .Q(ws2813_out_c_17)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_158), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_158), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_158), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n14081), .Z(n6954)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n14046), 
         .D(state[0]), .Z(sclk_c_enable_1530)) /* synthesis lut_function=(A (B)+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h9888;
    LUT4 i38462_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n14081), .Z(sclk_c_enable_158)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38462_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    L6MUX21 i37982 (.D0(n53184), .D1(n53185), .SD(bit_counter[2]), .Z(n53188));
    L6MUX21 i37983 (.D0(n53186), .D1(n53187), .SD(bit_counter[2]), .Z(n53189));
    LUT4 mux_2837_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n14081), .Z(n54968)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2837_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2837_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n14081), .Z(n54967)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2837_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 mux_2837_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14081), .Z(n54872)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2837_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2837_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14046), .Z(n54871)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2837_i3_4_lut_else_4_lut.init = 16'hd0f2;
    L6MUX21 i38155 (.D0(n53359), .D1(n53360), .SD(bit_counter[2]), .Z(n53361));
    LUT4 mux_2847_i2_4_lut (.A(n68), .B(n15113[0]), .C(n10392), .D(n52664), 
         .Z(n10393[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2847_i4_4_lut (.A(n37745), .B(n54696), .C(n10392), .D(n4), 
         .Z(n10393[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42686), .B(n54576), .C(n447[3]), .D(n54701), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2847_i8_4_lut (.A(n10217[7]), .B(n54696), .C(n10392), .D(n54576), 
         .Z(n10393[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i8_4_lut.init = 16'h303a;
    FD1P3IX pixel_i0 (.D(\Q[17] [0]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    LUT4 mux_2847_i9_4_lut (.A(n10217[8]), .B(n54696), .C(n10392), .D(n54576), 
         .Z(n10393[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i9_4_lut.init = 16'h303a;
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 mux_2847_i10_4_lut (.A(n76), .B(n54696), .C(n10392), .D(n54576), 
         .Z(n10393[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i10_4_lut.init = 16'h303a;
    LUT4 mux_2847_i13_4_lut (.A(n54576), .B(n54696), .C(n10392), .D(n103), 
         .Z(n10393[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i13_4_lut.init = 16'h3530;
    FD1P3AX delay_counter_i0_i1 (.D(n10393[1]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n10393[3]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n10393[7]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n10393[8]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n10393[9]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n10393[12]), .SP(sclk_c_enable_1745), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n42686), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_666 (.A(state[2]), .B(n42686), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_666.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_667 (.A(state[2]), .B(n42686), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_667.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_668 (.A(state[2]), .B(n42686), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_668.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_669 (.A(state[2]), .B(n42686), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_669.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_670 (.A(state[2]), .B(n42686), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_670.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_671 (.A(state[2]), .B(n42686), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_671.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_672 (.A(state[2]), .B(n42686), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_672.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_673 (.A(state[2]), .B(n42686), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_673.init = 16'h1010;
    LUT4 mux_2110_i2_4_lut_4_lut (.A(n54696), .B(n54701), .C(n6954), .D(n14046), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2110_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 i1_3_lut_4_lut (.A(n54565), .B(n54770), .C(n447[7]), .D(n54701), 
         .Z(n10217[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_674 (.A(n54565), .B(n54770), .C(n447[8]), 
         .D(n54701), .Z(n10217[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_674.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_675 (.A(n54565), .B(n54770), .C(n447[9]), 
         .D(n54701), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_675.init = 16'hf888;
    PFUMX i37978 (.BLUT(n53176), .ALUT(n53177), .C0(bit_counter[1]), .Z(n53184));
    LUT4 i38152_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38152_3_lut.init = 16'hcaca;
    PFUMX i37979 (.BLUT(n53178), .ALUT(n53179), .C0(bit_counter[1]), .Z(n53185));
    LUT4 i38151_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38151_3_lut.init = 16'hcaca;
    LUT4 i38150_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38150_3_lut.init = 16'hcaca;
    PFUMX i37980 (.BLUT(n53180), .ALUT(n53181), .C0(bit_counter[1]), .Z(n53186));
    LUT4 i38149_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38149_3_lut.init = 16'hcaca;
    PFUMX i37981 (.BLUT(n53182), .ALUT(n53183), .C0(bit_counter[1]), .Z(n53187));
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54636), .C(n14081), .D(n54770), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    FD1P3IX pixel_i23 (.D(\Q[17] [23]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[17] [22]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[17] [21]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[17] [20]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[17] [19]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[17] [18]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[17] [17]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[17] [16]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[17] [15]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54770), .B(state[1]), .C(n54636), .D(n54635), 
         .Z(n52664)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 i23959_2_lut_4_lut (.A(n54635), .B(state[0]), .C(state[1]), .D(n10392), 
         .Z(n36171)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23959_2_lut_4_lut.init = 16'hfd00;
    LUT4 i37977_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37977_3_lut.init = 16'hcaca;
    LUT4 i37976_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37976_3_lut.init = 16'hcaca;
    LUT4 i37975_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37975_3_lut.init = 16'hcaca;
    LUT4 i37974_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37974_3_lut.init = 16'hcaca;
    LUT4 i37973_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37973_3_lut.init = 16'hcaca;
    LUT4 i37972_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37972_3_lut.init = 16'hcaca;
    LUT4 i37971_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37971_3_lut.init = 16'hcaca;
    LUT4 i37970_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37970_3_lut.init = 16'hcaca;
    FD1P3IX pixel_i14 (.D(\Q[17] [14]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[17] [13]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[17] [12]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[17] [11]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[17] [10]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[17] [9]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[17] [8]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[17] [7]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[17] [6]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[17] [5]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[17] [4]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[17] [3]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[17] [2]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[17] [1]), .SP(sclk_c_enable_1563), .CD(n36353), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1530), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    L6MUX21 i37984 (.D0(n53188), .D1(n53189), .SD(bit_counter[3]), .Z(n53190));
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1563), 
            .CD(n36353), .CK(sclk_c), .Q(\RdAddress[17] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1594), .CD(n36353), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_912), .SP(sclk_c_enable_1594), .CD(n36353), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1594), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    PFUMX i38153 (.BLUT(n53355), .ALUT(n53356), .C0(bit_counter[1]), .Z(n53359));
    PFUMX i38154 (.BLUT(n53357), .ALUT(n53358), .C0(bit_counter[1]), .Z(n53360));
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1745), 
            .CD(n36175), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1745), .CD(n36175), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1745), .CD(n36175), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54969), .SP(sclk_c_enable_1745), .CD(n36171), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54873), .SP(sclk_c_enable_1745), .CD(n36171), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=322, LSE_RLINE=322 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i38426_2_lut_rep_747 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1594)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38426_2_lut_rep_747.init = 16'h9999;
    CCU2D add_3136_33 (.A0(bit_counter[31]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47935), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_33.INIT0 = 16'h5999;
    defparam add_3136_33.INIT1 = 16'h0000;
    defparam add_3136_33.INJECT1_0 = "NO";
    defparam add_3136_33.INJECT1_1 = "NO";
    CCU2D add_3136_31 (.A0(bit_counter[29]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47934), .COUT(n47935), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_31.INIT0 = 16'h5999;
    defparam add_3136_31.INIT1 = 16'h5999;
    defparam add_3136_31.INJECT1_0 = "NO";
    defparam add_3136_31.INJECT1_1 = "NO";
    CCU2D add_3136_29 (.A0(bit_counter[27]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47933), .COUT(n47934), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_29.INIT0 = 16'h5999;
    defparam add_3136_29.INIT1 = 16'h5999;
    defparam add_3136_29.INJECT1_0 = "NO";
    defparam add_3136_29.INJECT1_1 = "NO";
    CCU2D add_3136_27 (.A0(bit_counter[25]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47932), .COUT(n47933), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_27.INIT0 = 16'h5999;
    defparam add_3136_27.INIT1 = 16'h5999;
    defparam add_3136_27.INJECT1_0 = "NO";
    defparam add_3136_27.INJECT1_1 = "NO";
    CCU2D add_3136_25 (.A0(bit_counter[23]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47931), .COUT(n47932), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_25.INIT0 = 16'h5999;
    defparam add_3136_25.INIT1 = 16'h5999;
    defparam add_3136_25.INJECT1_0 = "NO";
    defparam add_3136_25.INJECT1_1 = "NO";
    CCU2D add_3136_23 (.A0(bit_counter[21]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47930), .COUT(n47931), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_23.INIT0 = 16'h5999;
    defparam add_3136_23.INIT1 = 16'h5999;
    defparam add_3136_23.INJECT1_0 = "NO";
    defparam add_3136_23.INJECT1_1 = "NO";
    CCU2D add_3136_21 (.A0(bit_counter[19]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47929), .COUT(n47930), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_21.INIT0 = 16'h5999;
    defparam add_3136_21.INIT1 = 16'h5999;
    defparam add_3136_21.INJECT1_0 = "NO";
    defparam add_3136_21.INJECT1_1 = "NO";
    CCU2D add_3136_19 (.A0(bit_counter[17]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47928), .COUT(n47929), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_19.INIT0 = 16'h5999;
    defparam add_3136_19.INIT1 = 16'h5999;
    defparam add_3136_19.INJECT1_0 = "NO";
    defparam add_3136_19.INJECT1_1 = "NO";
    CCU2D add_3136_17 (.A0(bit_counter[15]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47927), .COUT(n47928), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_17.INIT0 = 16'h5999;
    defparam add_3136_17.INIT1 = 16'h5999;
    defparam add_3136_17.INJECT1_0 = "NO";
    defparam add_3136_17.INJECT1_1 = "NO";
    LUT4 i25541_1_lut_rep_756 (.A(state[2]), .Z(n54759)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25541_1_lut_rep_756.init = 16'h5555;
    LUT4 i29990_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i29990_3_lut_3_lut.init = 16'h5151;
    CCU2D add_3136_15 (.A0(bit_counter[13]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47926), .COUT(n47927), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_15.INIT0 = 16'h5999;
    defparam add_3136_15.INIT1 = 16'h5999;
    defparam add_3136_15.INJECT1_0 = "NO";
    defparam add_3136_15.INJECT1_1 = "NO";
    CCU2D add_3136_13 (.A0(bit_counter[11]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47925), .COUT(n47926), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_13.INIT0 = 16'h5999;
    defparam add_3136_13.INIT1 = 16'h5999;
    defparam add_3136_13.INJECT1_0 = "NO";
    defparam add_3136_13.INJECT1_1 = "NO";
    CCU2D add_3136_11 (.A0(bit_counter[9]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47924), .COUT(n47925), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_11.INIT0 = 16'h5999;
    defparam add_3136_11.INIT1 = 16'h5999;
    defparam add_3136_11.INJECT1_0 = "NO";
    defparam add_3136_11.INJECT1_1 = "NO";
    CCU2D add_3136_9 (.A0(bit_counter[7]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47923), .COUT(n47924), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_9.INIT0 = 16'h5999;
    defparam add_3136_9.INIT1 = 16'h5999;
    defparam add_3136_9.INJECT1_0 = "NO";
    defparam add_3136_9.INJECT1_1 = "NO";
    CCU2D add_3136_7 (.A0(bit_counter[5]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47922), .COUT(n47923), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_7.INIT0 = 16'h5999;
    defparam add_3136_7.INIT1 = 16'h5999;
    defparam add_3136_7.INJECT1_0 = "NO";
    defparam add_3136_7.INJECT1_1 = "NO";
    CCU2D add_3136_5 (.A0(bit_counter[3]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47921), .COUT(n47922), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_5.INIT0 = 16'h5999;
    defparam add_3136_5.INIT1 = 16'h5999;
    defparam add_3136_5.INJECT1_0 = "NO";
    defparam add_3136_5.INJECT1_1 = "NO";
    CCU2D add_3136_3 (.A0(bit_counter[1]), .B0(n14046), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n14046), .C1(GND_net), 
          .D1(GND_net), .CIN(n47920), .COUT(n47921), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_3.INIT0 = 16'h5999;
    defparam add_3136_3.INIT1 = 16'h5999;
    defparam add_3136_3.INJECT1_0 = "NO";
    defparam add_3136_3.INJECT1_1 = "NO";
    CCU2D add_3136_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n14046), .C1(GND_net), .D1(GND_net), 
          .COUT(n47920), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3136_1.INIT0 = 16'hF000;
    defparam add_3136_1.INIT1 = 16'h5999;
    defparam add_3136_1.INJECT1_0 = "NO";
    defparam add_3136_1.INJECT1_1 = "NO";
    LUT4 i28790_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28790_2_lut.init = 16'hbbbb;
    LUT4 i28789_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_912)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28789_2_lut.init = 16'hbbbb;
    LUT4 mux_2847_i1_4_lut (.A(n69), .B(n15113[0]), .C(n10392), .D(n52664), 
         .Z(n10393[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2847_i1_4_lut.init = 16'hcfca;
    LUT4 i2859_3_lut (.A(state[2]), .B(state[1]), .C(n14081), .Z(n10392)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2859_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42686)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i107_3_lut_4_lut (.A(n42686), .B(n14046), .C(n54701), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 i23983_4_lut (.A(sclk_c_enable_1745), .B(n54701), .C(n10392), 
         .D(n54576), .Z(n36175)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23983_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_rep_698_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54701)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_698_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_676 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_676.init = 16'he0f0;
    LUT4 i1_2_lut_rep_767 (.A(state[2]), .B(state[0]), .Z(n54770)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_767.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_677 (.A(state[2]), .B(state[0]), .C(n14046), 
         .D(state[1]), .Z(n37745)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_677.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_adj_678 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_678.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_679 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_679.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_680 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_680.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_681 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_681.init = 16'h4040;
    PFUMX i38889 (.BLUT(n54871), .ALUT(n54872), .C0(state[1]), .Z(n54873));
    LUT4 i1_2_lut_3_lut_adj_682 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_682.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_683 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_683.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_684 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_684.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_685 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_685.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_686 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_686.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_687 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_687.init = 16'h4040;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_688 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_688.init = 16'h4040;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48083), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48082), .COUT(n48083), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_689 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_689.init = 16'h4040;
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48081), .COUT(n48082), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48080), .COUT(n48081), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_690 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_690.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_691 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_691.init = 16'h4040;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53190), .B(n53361), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_3_lut_adj_692 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_692.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_693 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_693.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_694 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_694.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_695 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_695.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_696 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_696.init = 16'h4040;
    LUT4 mux_2110_i1_4_lut (.A(n54636), .B(n54696), .C(n6954), .D(n54701), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2110_i1_4_lut.init = 16'h3f3a;
    LUT4 i1_2_lut_3_lut_adj_697 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_697.init = 16'h4040;
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48079), .COUT(n48080), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48078), .COUT(n48079), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48077), .COUT(n48078), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48076), .COUT(n48077), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_698 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_698.init = 16'h4040;
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48075), .COUT(n48076), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48074), .COUT(n48075), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48073), .COUT(n48074), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48072), .COUT(n48073), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_699 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_699.init = 16'h4040;
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48071), .COUT(n48072), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48070), .COUT(n48071), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_700 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_700.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_701 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_701.init = 16'h4040;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48069), .COUT(n48070), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_702 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_702.init = 16'h4040;
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48068), .COUT(n48069), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_703 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_703.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_704 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_704.init = 16'h4040;
    CCU2D add_33940_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48721), 
          .S0(n14081));
    defparam add_33940_cout.INIT0 = 16'h0000;
    defparam add_33940_cout.INIT1 = 16'h0000;
    defparam add_33940_cout.INJECT1_0 = "NO";
    defparam add_33940_cout.INJECT1_1 = "NO";
    CCU2D add_33940_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48720), .COUT(n48721));
    defparam add_33940_31.INIT0 = 16'hf555;
    defparam add_33940_31.INIT1 = 16'h5555;
    defparam add_33940_31.INJECT1_0 = "NO";
    defparam add_33940_31.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48068), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_33940_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48719), .COUT(n48720));
    defparam add_33940_29.INIT0 = 16'hf555;
    defparam add_33940_29.INIT1 = 16'hf555;
    defparam add_33940_29.INJECT1_0 = "NO";
    defparam add_33940_29.INJECT1_1 = "NO";
    CCU2D add_33940_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48718), .COUT(n48719));
    defparam add_33940_27.INIT0 = 16'hf555;
    defparam add_33940_27.INIT1 = 16'hf555;
    defparam add_33940_27.INJECT1_0 = "NO";
    defparam add_33940_27.INJECT1_1 = "NO";
    CCU2D add_33940_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48717), .COUT(n48718));
    defparam add_33940_25.INIT0 = 16'hf555;
    defparam add_33940_25.INIT1 = 16'hf555;
    defparam add_33940_25.INJECT1_0 = "NO";
    defparam add_33940_25.INJECT1_1 = "NO";
    CCU2D add_33940_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48716), .COUT(n48717));
    defparam add_33940_23.INIT0 = 16'hf555;
    defparam add_33940_23.INIT1 = 16'hf555;
    defparam add_33940_23.INJECT1_0 = "NO";
    defparam add_33940_23.INJECT1_1 = "NO";
    CCU2D add_33940_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48715), .COUT(n48716));
    defparam add_33940_21.INIT0 = 16'hf555;
    defparam add_33940_21.INIT1 = 16'hf555;
    defparam add_33940_21.INJECT1_0 = "NO";
    defparam add_33940_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_705 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_705.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_706 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_706.init = 16'h4040;
    CCU2D add_33940_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48714), .COUT(n48715));
    defparam add_33940_19.INIT0 = 16'hf555;
    defparam add_33940_19.INIT1 = 16'hf555;
    defparam add_33940_19.INJECT1_0 = "NO";
    defparam add_33940_19.INJECT1_1 = "NO";
    CCU2D add_33940_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48713), .COUT(n48714));
    defparam add_33940_17.INIT0 = 16'hf555;
    defparam add_33940_17.INIT1 = 16'hf555;
    defparam add_33940_17.INJECT1_0 = "NO";
    defparam add_33940_17.INJECT1_1 = "NO";
    CCU2D add_33940_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48712), .COUT(n48713));
    defparam add_33940_15.INIT0 = 16'hf555;
    defparam add_33940_15.INIT1 = 16'hf555;
    defparam add_33940_15.INJECT1_0 = "NO";
    defparam add_33940_15.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48066), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48065), .COUT(n48066), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_707 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_707.init = 16'h4040;
    CCU2D add_33940_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48711), .COUT(n48712));
    defparam add_33940_13.INIT0 = 16'hf555;
    defparam add_33940_13.INIT1 = 16'hf555;
    defparam add_33940_13.INJECT1_0 = "NO";
    defparam add_33940_13.INJECT1_1 = "NO";
    CCU2D add_33940_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48710), .COUT(n48711));
    defparam add_33940_11.INIT0 = 16'hf555;
    defparam add_33940_11.INIT1 = 16'hf555;
    defparam add_33940_11.INJECT1_0 = "NO";
    defparam add_33940_11.INJECT1_1 = "NO";
    CCU2D add_33940_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48709), .COUT(n48710));
    defparam add_33940_9.INIT0 = 16'hf555;
    defparam add_33940_9.INIT1 = 16'hf555;
    defparam add_33940_9.INJECT1_0 = "NO";
    defparam add_33940_9.INJECT1_1 = "NO";
    CCU2D add_33940_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48708), .COUT(n48709));
    defparam add_33940_7.INIT0 = 16'hf555;
    defparam add_33940_7.INIT1 = 16'hf555;
    defparam add_33940_7.INJECT1_0 = "NO";
    defparam add_33940_7.INJECT1_1 = "NO";
    CCU2D add_33940_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48707), .COUT(n48708));
    defparam add_33940_5.INIT0 = 16'hf555;
    defparam add_33940_5.INIT1 = 16'hf555;
    defparam add_33940_5.INJECT1_0 = "NO";
    defparam add_33940_5.INJECT1_1 = "NO";
    CCU2D add_33940_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48706), .COUT(n48707));
    defparam add_33940_3.INIT0 = 16'hf555;
    defparam add_33940_3.INIT1 = 16'hf555;
    defparam add_33940_3.INJECT1_0 = "NO";
    defparam add_33940_3.INJECT1_1 = "NO";
    CCU2D add_33940_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48706));
    defparam add_33940_1.INIT0 = 16'hF000;
    defparam add_33940_1.INIT1 = 16'ha666;
    defparam add_33940_1.INJECT1_0 = "NO";
    defparam add_33940_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_693_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54696)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_693_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_rep_688_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1563)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_688_4_lut_3_lut.init = 16'h8989;
    LUT4 i24204_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36353)) /* synthesis lut_function=(A (B)) */ ;
    defparam i24204_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_708 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15113[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_708.init = 16'h7070;
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48064), .COUT(n48065), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48063), .COUT(n48064), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48063), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n14081), 
         .Z(sclk_c_enable_155)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_rep_633 (.A(n42686), .B(n14046), .Z(n54636)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_633.init = 16'h8888;
    LUT4 i1_2_lut_rep_632 (.A(state[2]), .B(n14081), .Z(n54635)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_632.init = 16'h4444;
    LUT4 i1_2_lut_rep_562_3_lut (.A(n42686), .B(n14046), .C(state[1]), 
         .Z(n54565)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_562_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_573_3_lut (.A(state[2]), .B(n14081), .C(state[1]), 
         .Z(n54576)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_573_3_lut.init = 16'h4040;
    LUT4 i38576_3_lut_rep_574_4_lut (.A(state[2]), .B(n14081), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1745)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38576_3_lut_rep_574_4_lut.init = 16'hfffb;
    PFUMX i38953 (.BLUT(n54967), .ALUT(n54968), .C0(state[0]), .Z(n54969));
    CCU2D add_33896_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48625), 
          .S0(n14046));
    defparam add_33896_cout.INIT0 = 16'h0000;
    defparam add_33896_cout.INIT1 = 16'h0000;
    defparam add_33896_cout.INJECT1_0 = "NO";
    defparam add_33896_cout.INJECT1_1 = "NO";
    CCU2D add_33896_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48624), .COUT(n48625));
    defparam add_33896_31.INIT0 = 16'hf555;
    defparam add_33896_31.INIT1 = 16'h5555;
    defparam add_33896_31.INJECT1_0 = "NO";
    defparam add_33896_31.INJECT1_1 = "NO";
    CCU2D add_33896_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48623), .COUT(n48624));
    defparam add_33896_29.INIT0 = 16'hf555;
    defparam add_33896_29.INIT1 = 16'hf555;
    defparam add_33896_29.INJECT1_0 = "NO";
    defparam add_33896_29.INJECT1_1 = "NO";
    CCU2D add_33896_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48622), .COUT(n48623));
    defparam add_33896_27.INIT0 = 16'hf555;
    defparam add_33896_27.INIT1 = 16'hf555;
    defparam add_33896_27.INJECT1_0 = "NO";
    defparam add_33896_27.INJECT1_1 = "NO";
    CCU2D add_33896_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48621), .COUT(n48622));
    defparam add_33896_25.INIT0 = 16'hf555;
    defparam add_33896_25.INIT1 = 16'hf555;
    defparam add_33896_25.INJECT1_0 = "NO";
    defparam add_33896_25.INJECT1_1 = "NO";
    CCU2D add_33896_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48620), .COUT(n48621));
    defparam add_33896_23.INIT0 = 16'hf555;
    defparam add_33896_23.INIT1 = 16'hf555;
    defparam add_33896_23.INJECT1_0 = "NO";
    defparam add_33896_23.INJECT1_1 = "NO";
    CCU2D add_33896_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48619), .COUT(n48620));
    defparam add_33896_21.INIT0 = 16'hf555;
    defparam add_33896_21.INIT1 = 16'hf555;
    defparam add_33896_21.INJECT1_0 = "NO";
    defparam add_33896_21.INJECT1_1 = "NO";
    CCU2D add_33896_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48618), .COUT(n48619));
    defparam add_33896_19.INIT0 = 16'hf555;
    defparam add_33896_19.INIT1 = 16'hf555;
    defparam add_33896_19.INJECT1_0 = "NO";
    defparam add_33896_19.INJECT1_1 = "NO";
    CCU2D add_33896_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48617), .COUT(n48618));
    defparam add_33896_17.INIT0 = 16'hf555;
    defparam add_33896_17.INIT1 = 16'hf555;
    defparam add_33896_17.INJECT1_0 = "NO";
    defparam add_33896_17.INJECT1_1 = "NO";
    CCU2D add_33896_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48616), .COUT(n48617));
    defparam add_33896_15.INIT0 = 16'hf555;
    defparam add_33896_15.INIT1 = 16'hf555;
    defparam add_33896_15.INJECT1_0 = "NO";
    defparam add_33896_15.INJECT1_1 = "NO";
    CCU2D add_33896_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48615), .COUT(n48616));
    defparam add_33896_13.INIT0 = 16'hf555;
    defparam add_33896_13.INIT1 = 16'hf555;
    defparam add_33896_13.INJECT1_0 = "NO";
    defparam add_33896_13.INJECT1_1 = "NO";
    CCU2D add_33896_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48614), .COUT(n48615));
    defparam add_33896_11.INIT0 = 16'hf555;
    defparam add_33896_11.INIT1 = 16'hf555;
    defparam add_33896_11.INJECT1_0 = "NO";
    defparam add_33896_11.INJECT1_1 = "NO";
    CCU2D add_33896_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48613), .COUT(n48614));
    defparam add_33896_9.INIT0 = 16'hf555;
    defparam add_33896_9.INIT1 = 16'hf555;
    defparam add_33896_9.INJECT1_0 = "NO";
    defparam add_33896_9.INJECT1_1 = "NO";
    CCU2D add_33896_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48612), .COUT(n48613));
    defparam add_33896_7.INIT0 = 16'hf555;
    defparam add_33896_7.INIT1 = 16'hf555;
    defparam add_33896_7.INJECT1_0 = "NO";
    defparam add_33896_7.INJECT1_1 = "NO";
    CCU2D add_33896_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48611), .COUT(n48612));
    defparam add_33896_5.INIT0 = 16'hf555;
    defparam add_33896_5.INIT1 = 16'hf555;
    defparam add_33896_5.INJECT1_0 = "NO";
    defparam add_33896_5.INJECT1_1 = "NO";
    CCU2D add_33896_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48610), .COUT(n48611));
    defparam add_33896_3.INIT0 = 16'hf555;
    defparam add_33896_3.INIT1 = 16'hf555;
    defparam add_33896_3.INJECT1_0 = "NO";
    defparam add_33896_3.INJECT1_1 = "NO";
    CCU2D add_33896_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48610));
    defparam add_33896_1.INIT0 = 16'hF000;
    defparam add_33896_1.INIT1 = 16'ha666;
    defparam add_33896_1.INJECT1_0 = "NO";
    defparam add_33896_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U26 
//

module \WS2812(48000000,"111111111")_U26  (sclk_c, \port_status[2] , ws2813_out_c_2, 
            GND_net, \Q[2] , \RdAddress[2] );
    input sclk_c;
    output \port_status[2] ;
    output ws2813_out_c_2;
    input GND_net;
    input [23:0]\Q[2] ;
    output [8:0]\RdAddress[2] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n52957, n52958;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n52962;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_873;
    wire [31:0]n7678;
    
    wire sclk_c_enable_27, n54784, sclk_c_enable_28, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_32;
    wire [2:0]state_2__N_104;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n47587;
    wire [31:0]n447;
    
    wire n47588, n47586, n47585, n47584, n47583, n47582, n42596, 
        n12996, n55530, n47581, n54916, n13031, n54905, n54904, 
        n27;
    wire [6:0]n15031;
    
    wire n54677, n52676, n54914, n54913, n54917, n15;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire n14, serial_N_437, n54953, n54952, n54987, n54986, n53254, 
        n53255, n53256, sclk_c_enable_1226, n52956, n52955, sclk_c_enable_1225, 
        n54837, sclk_c_enable_1224;
    wire [8:0]cur_pixel_8__N_107;
    wire [31:0]bit_counter_31__N_172;
    
    wire n1, n1_adj_911, n34750, n34746, n54915, n54906, n52954, 
        n52959, n52960, n52963, n52961, n52964, n52953, n54856, 
        n54857, n54618, n54735;
    wire [31:0]n7502;
    
    wire n52952, n52951, n54736, n29;
    wire [8:0]n118;
    
    wire n42552;
    wire [31:0]bit_counter_31__N_204;
    
    wire n47580, n47579, n47578, n47577, n53253, n53252, n53251, 
        n53250, n47575, n47574, n47573, n47572, n48242, n48241, 
        n48240, n48239, n48238, n48237, n48236, n48235, n48234, 
        n48233, n48232, n48231, n48230, n48229, n48228, n48227, 
        n52965, n48849, n48848, n48847, n48846, n48845, n48844, 
        n48843, n48842, n48841, n48840, n48839, n48838, n48837, 
        n48836, n48835, n48834, n48785, n48784, n48783, n48782, 
        n48781, n48780, n48779, n48778, n48777, n48776, n48775, 
        n48774, n48773, n48772, n48771, n48770, n47592, n47591, 
        n47590, n47589;
    
    PFUMX i37756 (.BLUT(n52957), .ALUT(n52958), .C0(bit_counter[1]), .Z(n52962));
    FD1P3AX delay_counter_i0_i0 (.D(n7678[0]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54784), .SP(sclk_c_enable_27), .CK(sclk_c), 
            .Q(\port_status[2] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_28), .CK(sclk_c), 
            .Q(ws2813_out_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_32), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_32), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_32), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i37752_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n52958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37752_3_lut.init = 16'hcaca;
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47587), .COUT(n47588), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47586), .COUT(n47587), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47585), .COUT(n47586), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47584), .COUT(n47585), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47583), .COUT(n47584), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47582), .COUT(n47583), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    LUT4 i29267_2_lut_rep_841 (.A(n42596), .B(n12996), .Z(n55530)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29267_2_lut_rep_841.init = 16'h8888;
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47581), .COUT(n47582), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut_else_2_lut_4_lut (.A(n42596), .B(n12996), 
         .C(state[0]), .D(state[2]), .Z(n54916)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_else_2_lut_4_lut.init = 16'h0070;
    LUT4 mux_2240_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13031), .Z(n54905)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2240_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2240_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n12996), .Z(n54904)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2240_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 mux_2250_i1_4_lut (.A(n27), .B(n15031[0]), .C(n54677), .D(n52676), 
         .Z(n7678[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i1_4_lut.init = 16'hcfca;
    LUT4 mux_2240_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13031), .Z(n54914)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam mux_2240_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2240_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13031), .Z(n54913)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam mux_2240_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 i1_3_lut_4_lut_4_lut_then_2_lut (.A(n13031), .B(state[2]), .Z(n54917)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_3_lut_4_lut_4_lut_then_2_lut.init = 16'h2222;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[7]), .C(n14), .D(cur_pixel[4]), 
         .Z(n42596)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i27502_1_lut_rep_781 (.A(state[2]), .Z(n54784)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27502_1_lut_rep_781.init = 16'h5555;
    LUT4 i28827_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28827_3_lut_3_lut.init = 16'h5151;
    LUT4 i6_4_lut (.A(cur_pixel[2]), .B(cur_pixel[8]), .C(cur_pixel[6]), 
         .D(cur_pixel[5]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[3]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 mux_2935_i3_then_3_lut (.A(state[2]), .B(state[0]), .C(n13031), 
         .Z(n54953)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam mux_2935_i3_then_3_lut.init = 16'h4040;
    LUT4 mux_2935_i3_else_3_lut (.A(state[2]), .B(state[0]), .C(n42596), 
         .D(n12996), .Z(n54952)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam mux_2935_i3_else_3_lut.init = 16'h4000;
    LUT4 mux_2935_i2_3_lut_4_lut_then_3_lut (.A(state[1]), .B(state[2]), 
         .C(n12996), .Z(n54987)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam mux_2935_i2_3_lut_4_lut_then_3_lut.init = 16'h0101;
    LUT4 mux_2935_i2_3_lut_4_lut_else_3_lut (.A(state[1]), .B(state[2]), 
         .C(n13031), .Z(n54986)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam mux_2935_i2_3_lut_4_lut_else_3_lut.init = 16'h2020;
    L6MUX21 i38050 (.D0(n53254), .D1(n53255), .SD(bit_counter[2]), .Z(n53256));
    LUT4 i38420_2_lut_rep_794 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1226)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38420_2_lut_rep_794.init = 16'h9999;
    LUT4 i37750_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n52956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37750_3_lut.init = 16'hcaca;
    LUT4 i37749_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n52955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37749_3_lut.init = 16'hcaca;
    FD1P3IX pixel_i23 (.D(\Q[2] [23]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[2] [22]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[2] [21]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[2] [20]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[2] [19]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[2] [18]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[2] [17]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[2] [16]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[2] [15]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[2] [14]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[2] [13]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[2] [12]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[2] [11]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[2] [10]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[2] [9]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[2] [8]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[2] [7]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[2] [6]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[2] [5]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[2] [4]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[2] [3]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[2] [2]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[2] [1]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1226), .CD(n54837), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_911), .SP(sclk_c_enable_1226), .CD(n54837), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_873), 
            .CD(n34750), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_873), .CD(n34750), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_873), .CD(n34750), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54915), .SP(sclk_c_enable_873), .CD(n34746), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54906), .SP(sclk_c_enable_873), .CD(n34746), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i1 (.D(n7678[1]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n7678[3]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n7678[7]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n7678[8]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n7678[9]), .SP(sclk_c_enable_873), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n7678[12]), .SP(sclk_c_enable_873), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i37748_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37748_3_lut.init = 16'hcaca;
    L6MUX21 i37757 (.D0(n52959), .D1(n52960), .SD(bit_counter[2]), .Z(n52963));
    L6MUX21 i37758 (.D0(n52961), .D1(n52962), .SD(bit_counter[2]), .Z(n52964));
    LUT4 i37747_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37747_3_lut.init = 16'hcaca;
    PFUMX i38879 (.BLUT(n54856), .ALUT(n54857), .C0(n55530), .Z(state_2__N_104[0]));
    LUT4 i1_2_lut_rep_615_3_lut (.A(state[2]), .B(n13031), .C(state[1]), 
         .Z(n54618)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_615_3_lut.init = 16'h4040;
    LUT4 mux_2234_i8_3_lut_4_lut (.A(n42596), .B(n12996), .C(n54735), 
         .D(n447[7]), .Z(n7502[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2234_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2234_i9_3_lut_4_lut (.A(n42596), .B(n12996), .C(n54735), 
         .D(n447[8]), .Z(n7502[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2234_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2234_i10_3_lut_4_lut (.A(n42596), .B(n12996), .C(n54735), 
         .D(n447[9]), .Z(n7502[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2234_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2234_i13_3_lut_4_lut (.A(n42596), .B(n12996), .C(n54735), 
         .D(n447[12]), .Z(n7502[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2234_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i2262_3_lut_rep_674 (.A(state[2]), .B(state[1]), .C(n13031), 
         .Z(n54677)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2262_3_lut_rep_674.init = 16'ha8a8;
    LUT4 i37746_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37746_3_lut.init = 16'hcaca;
    LUT4 i37745_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37745_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n27)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i2_2_lut_rep_733_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54736)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2_2_lut_rep_733_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_627 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n29)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_627.init = 16'he0f0;
    LUT4 i38630_2_lut_rep_552_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(n13031), .D(state[2]), .Z(sclk_c_enable_873)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i38630_2_lut_rep_552_2_lut_3_lut_4_lut.init = 16'hffef;
    LUT4 i22534_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut (.A(state[1]), .B(n13031), 
         .C(state[2]), .Z(n34746)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i22534_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut.init = 16'he0e0;
    FD1P3IX pixel_i0 (.D(\Q[2] [0]), .SP(sclk_c_enable_1225), .CD(n54837), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1224), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1225), 
            .CD(n54837), .CK(sclk_c), .Q(\RdAddress[2] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1226), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=157, LSE_RLINE=157 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i27508_3_lut_3_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(sclk_c_enable_1225)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam i27508_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n42596), .C(n118[8]), .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_628 (.A(state[2]), .B(n42596), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_628.init = 16'h1010;
    LUT4 i1_2_lut_rep_834 (.A(state[2]), .B(state[1]), .Z(n54837)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_834.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_629 (.A(state[2]), .B(n42596), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_629.init = 16'h1010;
    LUT4 i30381_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42552)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i30381_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_adj_630 (.A(state[2]), .B(n42596), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_630.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_631 (.A(state[2]), .B(n42596), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_631.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_632 (.A(state[2]), .B(n42596), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_632.init = 16'h1010;
    LUT4 i28692_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15031[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28692_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13031), 
         .Z(sclk_c_enable_28)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_3_lut_adj_633 (.A(state[2]), .B(n42596), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_633.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_634 (.A(state[2]), .B(n42596), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_634.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_635 (.A(state[2]), .B(n42596), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_635.init = 16'h1010;
    LUT4 i37683_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13031), 
         .D(state[1]), .Z(sclk_c_enable_32)) /* synthesis lut_function=(A (C+(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i37683_3_lut_4_lut_4_lut_4_lut.init = 16'hfaf4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n12996), 
         .D(state[1]), .Z(sclk_c_enable_1224)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_rep_732_3_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .Z(n54735)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_732_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_3_lut_adj_636 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_636.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_637 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_637.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_638 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_638.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_639 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_639.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_640 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_640.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_641 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_641.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_642 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_642.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_643 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_643.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_644 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_644.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_645 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_645.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_646 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_646.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_647 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_647.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_648 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_648.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_649 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_649.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_650 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_650.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_651 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_651.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_652 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_652.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_653 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_653.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_654 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_654.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_655 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_655.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_656 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_656.init = 16'h4040;
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47580), .COUT(n47581), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_657 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_657.init = 16'h4040;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47579), .COUT(n47580), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_658 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_658.init = 16'h4040;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47578), .COUT(n47579), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_659 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_659.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_660 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_660.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_661 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_661.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_662 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_662.init = 16'h4040;
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47577), .COUT(n47578), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_663 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_663.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_664 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_664.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_665 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_665.init = 16'h4040;
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47577), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i38047_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38047_3_lut.init = 16'hcaca;
    LUT4 i38046_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38046_3_lut.init = 16'hcaca;
    LUT4 i38045_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38045_3_lut.init = 16'hcaca;
    LUT4 i38044_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38044_3_lut.init = 16'hcaca;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47575), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47574), .COUT(n47575), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    PFUMX i38048 (.BLUT(n53250), .ALUT(n53251), .C0(bit_counter[1]), .Z(n53254));
    PFUMX i38049 (.BLUT(n53252), .ALUT(n53253), .C0(bit_counter[1]), .Z(n53255));
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47573), .COUT(n47574), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47572), .COUT(n47573), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47572), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3106_33 (.A0(bit_counter[31]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48242), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_33.INIT0 = 16'h5999;
    defparam add_3106_33.INIT1 = 16'h0000;
    defparam add_3106_33.INJECT1_0 = "NO";
    defparam add_3106_33.INJECT1_1 = "NO";
    CCU2D add_3106_31 (.A0(bit_counter[29]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48241), .COUT(n48242), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_31.INIT0 = 16'h5999;
    defparam add_3106_31.INIT1 = 16'h5999;
    defparam add_3106_31.INJECT1_0 = "NO";
    defparam add_3106_31.INJECT1_1 = "NO";
    CCU2D add_3106_29 (.A0(bit_counter[27]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48240), .COUT(n48241), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_29.INIT0 = 16'h5999;
    defparam add_3106_29.INIT1 = 16'h5999;
    defparam add_3106_29.INJECT1_0 = "NO";
    defparam add_3106_29.INJECT1_1 = "NO";
    CCU2D add_3106_27 (.A0(bit_counter[25]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48239), .COUT(n48240), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_27.INIT0 = 16'h5999;
    defparam add_3106_27.INIT1 = 16'h5999;
    defparam add_3106_27.INJECT1_0 = "NO";
    defparam add_3106_27.INJECT1_1 = "NO";
    CCU2D add_3106_25 (.A0(bit_counter[23]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48238), .COUT(n48239), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_25.INIT0 = 16'h5999;
    defparam add_3106_25.INIT1 = 16'h5999;
    defparam add_3106_25.INJECT1_0 = "NO";
    defparam add_3106_25.INJECT1_1 = "NO";
    CCU2D add_3106_23 (.A0(bit_counter[21]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48237), .COUT(n48238), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_23.INIT0 = 16'h5999;
    defparam add_3106_23.INIT1 = 16'h5999;
    defparam add_3106_23.INJECT1_0 = "NO";
    defparam add_3106_23.INJECT1_1 = "NO";
    CCU2D add_3106_21 (.A0(bit_counter[19]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48236), .COUT(n48237), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_21.INIT0 = 16'h5999;
    defparam add_3106_21.INIT1 = 16'h5999;
    defparam add_3106_21.INJECT1_0 = "NO";
    defparam add_3106_21.INJECT1_1 = "NO";
    CCU2D add_3106_19 (.A0(bit_counter[17]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48235), .COUT(n48236), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_19.INIT0 = 16'h5999;
    defparam add_3106_19.INIT1 = 16'h5999;
    defparam add_3106_19.INJECT1_0 = "NO";
    defparam add_3106_19.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    CCU2D add_3106_17 (.A0(bit_counter[15]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48234), .COUT(n48235), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_17.INIT0 = 16'h5999;
    defparam add_3106_17.INIT1 = 16'h5999;
    defparam add_3106_17.INJECT1_0 = "NO";
    defparam add_3106_17.INJECT1_1 = "NO";
    CCU2D add_3106_15 (.A0(bit_counter[13]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48233), .COUT(n48234), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_15.INIT0 = 16'h5999;
    defparam add_3106_15.INIT1 = 16'h5999;
    defparam add_3106_15.INJECT1_0 = "NO";
    defparam add_3106_15.INJECT1_1 = "NO";
    CCU2D add_3106_13 (.A0(bit_counter[11]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48232), .COUT(n48233), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_13.INIT0 = 16'h5999;
    defparam add_3106_13.INIT1 = 16'h5999;
    defparam add_3106_13.INJECT1_0 = "NO";
    defparam add_3106_13.INJECT1_1 = "NO";
    CCU2D add_3106_11 (.A0(bit_counter[9]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48231), .COUT(n48232), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_11.INIT0 = 16'h5999;
    defparam add_3106_11.INIT1 = 16'h5999;
    defparam add_3106_11.INJECT1_0 = "NO";
    defparam add_3106_11.INJECT1_1 = "NO";
    CCU2D add_3106_9 (.A0(bit_counter[7]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48230), .COUT(n48231), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_9.INIT0 = 16'h5999;
    defparam add_3106_9.INIT1 = 16'h5999;
    defparam add_3106_9.INJECT1_0 = "NO";
    defparam add_3106_9.INJECT1_1 = "NO";
    CCU2D add_3106_7 (.A0(bit_counter[5]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48229), .COUT(n48230), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_7.INIT0 = 16'h5999;
    defparam add_3106_7.INIT1 = 16'h5999;
    defparam add_3106_7.INJECT1_0 = "NO";
    defparam add_3106_7.INJECT1_1 = "NO";
    CCU2D add_3106_5 (.A0(bit_counter[3]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48228), .COUT(n48229), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_5.INIT0 = 16'h5999;
    defparam add_3106_5.INIT1 = 16'h5999;
    defparam add_3106_5.INJECT1_0 = "NO";
    defparam add_3106_5.INJECT1_1 = "NO";
    CCU2D add_3106_3 (.A0(bit_counter[1]), .B0(n12996), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n12996), .C1(GND_net), 
          .D1(GND_net), .CIN(n48227), .COUT(n48228), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_3.INIT0 = 16'h5999;
    defparam add_3106_3.INIT1 = 16'h5999;
    defparam add_3106_3.INJECT1_0 = "NO";
    defparam add_3106_3.INJECT1_1 = "NO";
    CCU2D add_3106_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n12996), .C1(GND_net), .D1(GND_net), 
          .COUT(n48227), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3106_1.INIT0 = 16'hF000;
    defparam add_3106_1.INIT1 = 16'h5999;
    defparam add_3106_1.INJECT1_0 = "NO";
    defparam add_3106_1.INJECT1_1 = "NO";
    LUT4 i28756_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28756_2_lut.init = 16'hbbbb;
    LUT4 i28757_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_911)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28757_2_lut.init = 16'hbbbb;
    L6MUX21 i37759 (.D0(n52963), .D1(n52964), .SD(bit_counter[3]), .Z(n52965));
    PFUMX i37753 (.BLUT(n52951), .ALUT(n52952), .C0(bit_counter[1]), .Z(n52959));
    LUT4 i22558_4_lut (.A(sclk_c_enable_873), .B(n54618), .C(n54677), 
         .D(n54735), .Z(n34750)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22558_4_lut.init = 16'haaa8;
    LUT4 mux_2935_i1_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(n13031), .Z(n54857)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B (C (D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2935_i1_4_lut_then_4_lut.init = 16'h175f;
    LUT4 mux_2935_i1_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(n13031), .Z(n54856)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B ((D)+!C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2935_i1_4_lut_else_4_lut.init = 16'h135b;
    LUT4 mux_2250_i2_4_lut (.A(n29), .B(n15031[0]), .C(n54677), .D(n52676), 
         .Z(n7678[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2250_i4_4_lut (.A(n7502[3]), .B(n42552), .C(n54677), .D(n54618), 
         .Z(n7678[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i4_4_lut.init = 16'h3f3a;
    LUT4 i29527_4_lut (.A(n42596), .B(n447[3]), .C(n54736), .D(n12996), 
         .Z(n7502[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29527_4_lut.init = 16'hcacf;
    LUT4 mux_2250_i8_4_lut (.A(n7502[7]), .B(n42552), .C(n54677), .D(n54618), 
         .Z(n7678[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i8_4_lut.init = 16'h303a;
    LUT4 mux_2250_i9_4_lut (.A(n7502[8]), .B(n42552), .C(n54677), .D(n54618), 
         .Z(n7678[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i9_4_lut.init = 16'h303a;
    LUT4 mux_2250_i10_4_lut (.A(n7502[9]), .B(n42552), .C(n54677), .D(n54618), 
         .Z(n7678[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i10_4_lut.init = 16'h303a;
    LUT4 mux_2250_i13_4_lut (.A(n7502[12]), .B(n42552), .C(n54677), .D(n54618), 
         .Z(n7678[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2250_i13_4_lut.init = 16'h303a;
    PFUMX i37754 (.BLUT(n52953), .ALUT(n52954), .C0(bit_counter[1]), .Z(n52960));
    CCU2D add_33935_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48849), 
          .S0(n13031));
    defparam add_33935_cout.INIT0 = 16'h0000;
    defparam add_33935_cout.INIT1 = 16'h0000;
    defparam add_33935_cout.INJECT1_0 = "NO";
    defparam add_33935_cout.INJECT1_1 = "NO";
    CCU2D add_33935_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48848), .COUT(n48849));
    defparam add_33935_31.INIT0 = 16'hf555;
    defparam add_33935_31.INIT1 = 16'h5555;
    defparam add_33935_31.INJECT1_0 = "NO";
    defparam add_33935_31.INJECT1_1 = "NO";
    CCU2D add_33935_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48847), .COUT(n48848));
    defparam add_33935_29.INIT0 = 16'hf555;
    defparam add_33935_29.INIT1 = 16'hf555;
    defparam add_33935_29.INJECT1_0 = "NO";
    defparam add_33935_29.INJECT1_1 = "NO";
    CCU2D add_33935_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48846), .COUT(n48847));
    defparam add_33935_27.INIT0 = 16'hf555;
    defparam add_33935_27.INIT1 = 16'hf555;
    defparam add_33935_27.INJECT1_0 = "NO";
    defparam add_33935_27.INJECT1_1 = "NO";
    CCU2D add_33935_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48845), .COUT(n48846));
    defparam add_33935_25.INIT0 = 16'hf555;
    defparam add_33935_25.INIT1 = 16'hf555;
    defparam add_33935_25.INJECT1_0 = "NO";
    defparam add_33935_25.INJECT1_1 = "NO";
    CCU2D add_33935_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48844), .COUT(n48845));
    defparam add_33935_23.INIT0 = 16'hf555;
    defparam add_33935_23.INIT1 = 16'hf555;
    defparam add_33935_23.INJECT1_0 = "NO";
    defparam add_33935_23.INJECT1_1 = "NO";
    CCU2D add_33935_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48843), .COUT(n48844));
    defparam add_33935_21.INIT0 = 16'hf555;
    defparam add_33935_21.INIT1 = 16'hf555;
    defparam add_33935_21.INJECT1_0 = "NO";
    defparam add_33935_21.INJECT1_1 = "NO";
    CCU2D add_33935_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48842), .COUT(n48843));
    defparam add_33935_19.INIT0 = 16'hf555;
    defparam add_33935_19.INIT1 = 16'hf555;
    defparam add_33935_19.INJECT1_0 = "NO";
    defparam add_33935_19.INJECT1_1 = "NO";
    CCU2D add_33935_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48841), .COUT(n48842));
    defparam add_33935_17.INIT0 = 16'hf555;
    defparam add_33935_17.INIT1 = 16'hf555;
    defparam add_33935_17.INJECT1_0 = "NO";
    defparam add_33935_17.INJECT1_1 = "NO";
    CCU2D add_33935_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48840), .COUT(n48841));
    defparam add_33935_15.INIT0 = 16'hf555;
    defparam add_33935_15.INIT1 = 16'hf555;
    defparam add_33935_15.INJECT1_0 = "NO";
    defparam add_33935_15.INJECT1_1 = "NO";
    CCU2D add_33935_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48839), .COUT(n48840));
    defparam add_33935_13.INIT0 = 16'hf555;
    defparam add_33935_13.INIT1 = 16'hf555;
    defparam add_33935_13.INJECT1_0 = "NO";
    defparam add_33935_13.INJECT1_1 = "NO";
    CCU2D add_33935_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48838), .COUT(n48839));
    defparam add_33935_11.INIT0 = 16'hf555;
    defparam add_33935_11.INIT1 = 16'hf555;
    defparam add_33935_11.INJECT1_0 = "NO";
    defparam add_33935_11.INJECT1_1 = "NO";
    CCU2D add_33935_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48837), .COUT(n48838));
    defparam add_33935_9.INIT0 = 16'hf555;
    defparam add_33935_9.INIT1 = 16'hf555;
    defparam add_33935_9.INJECT1_0 = "NO";
    defparam add_33935_9.INJECT1_1 = "NO";
    CCU2D add_33935_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48836), .COUT(n48837));
    defparam add_33935_7.INIT0 = 16'hf555;
    defparam add_33935_7.INIT1 = 16'hf555;
    defparam add_33935_7.INJECT1_0 = "NO";
    defparam add_33935_7.INJECT1_1 = "NO";
    CCU2D add_33935_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48835), .COUT(n48836));
    defparam add_33935_5.INIT0 = 16'hf555;
    defparam add_33935_5.INIT1 = 16'hf555;
    defparam add_33935_5.INJECT1_0 = "NO";
    defparam add_33935_5.INJECT1_1 = "NO";
    CCU2D add_33935_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48834), .COUT(n48835));
    defparam add_33935_3.INIT0 = 16'hf555;
    defparam add_33935_3.INIT1 = 16'hf555;
    defparam add_33935_3.INJECT1_0 = "NO";
    defparam add_33935_3.INJECT1_1 = "NO";
    CCU2D add_33935_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48834));
    defparam add_33935_1.INIT0 = 16'hF000;
    defparam add_33935_1.INIT1 = 16'ha666;
    defparam add_33935_1.INJECT1_0 = "NO";
    defparam add_33935_1.INJECT1_1 = "NO";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n52965), .B(n53256), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    CCU2D add_33937_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48785), 
          .S0(n12996));
    defparam add_33937_cout.INIT0 = 16'h0000;
    defparam add_33937_cout.INIT1 = 16'h0000;
    defparam add_33937_cout.INJECT1_0 = "NO";
    defparam add_33937_cout.INJECT1_1 = "NO";
    CCU2D add_33937_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48784), .COUT(n48785));
    defparam add_33937_31.INIT0 = 16'hf555;
    defparam add_33937_31.INIT1 = 16'h5555;
    defparam add_33937_31.INJECT1_0 = "NO";
    defparam add_33937_31.INJECT1_1 = "NO";
    CCU2D add_33937_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48783), .COUT(n48784));
    defparam add_33937_29.INIT0 = 16'hf555;
    defparam add_33937_29.INIT1 = 16'hf555;
    defparam add_33937_29.INJECT1_0 = "NO";
    defparam add_33937_29.INJECT1_1 = "NO";
    CCU2D add_33937_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48782), .COUT(n48783));
    defparam add_33937_27.INIT0 = 16'hf555;
    defparam add_33937_27.INIT1 = 16'hf555;
    defparam add_33937_27.INJECT1_0 = "NO";
    defparam add_33937_27.INJECT1_1 = "NO";
    CCU2D add_33937_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48781), .COUT(n48782));
    defparam add_33937_25.INIT0 = 16'hf555;
    defparam add_33937_25.INIT1 = 16'hf555;
    defparam add_33937_25.INJECT1_0 = "NO";
    defparam add_33937_25.INJECT1_1 = "NO";
    CCU2D add_33937_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48780), .COUT(n48781));
    defparam add_33937_23.INIT0 = 16'hf555;
    defparam add_33937_23.INIT1 = 16'hf555;
    defparam add_33937_23.INJECT1_0 = "NO";
    defparam add_33937_23.INJECT1_1 = "NO";
    CCU2D add_33937_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48779), .COUT(n48780));
    defparam add_33937_21.INIT0 = 16'hf555;
    defparam add_33937_21.INIT1 = 16'hf555;
    defparam add_33937_21.INJECT1_0 = "NO";
    defparam add_33937_21.INJECT1_1 = "NO";
    CCU2D add_33937_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48778), .COUT(n48779));
    defparam add_33937_19.INIT0 = 16'hf555;
    defparam add_33937_19.INIT1 = 16'hf555;
    defparam add_33937_19.INJECT1_0 = "NO";
    defparam add_33937_19.INJECT1_1 = "NO";
    CCU2D add_33937_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48777), .COUT(n48778));
    defparam add_33937_17.INIT0 = 16'hf555;
    defparam add_33937_17.INIT1 = 16'hf555;
    defparam add_33937_17.INJECT1_0 = "NO";
    defparam add_33937_17.INJECT1_1 = "NO";
    CCU2D add_33937_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48776), .COUT(n48777));
    defparam add_33937_15.INIT0 = 16'hf555;
    defparam add_33937_15.INIT1 = 16'hf555;
    defparam add_33937_15.INJECT1_0 = "NO";
    defparam add_33937_15.INJECT1_1 = "NO";
    CCU2D add_33937_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48775), .COUT(n48776));
    defparam add_33937_13.INIT0 = 16'hf555;
    defparam add_33937_13.INIT1 = 16'hf555;
    defparam add_33937_13.INJECT1_0 = "NO";
    defparam add_33937_13.INJECT1_1 = "NO";
    CCU2D add_33937_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48774), .COUT(n48775));
    defparam add_33937_11.INIT0 = 16'hf555;
    defparam add_33937_11.INIT1 = 16'hf555;
    defparam add_33937_11.INJECT1_0 = "NO";
    defparam add_33937_11.INJECT1_1 = "NO";
    CCU2D add_33937_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48773), .COUT(n48774));
    defparam add_33937_9.INIT0 = 16'hf555;
    defparam add_33937_9.INIT1 = 16'hf555;
    defparam add_33937_9.INJECT1_0 = "NO";
    defparam add_33937_9.INJECT1_1 = "NO";
    CCU2D add_33937_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48772), .COUT(n48773));
    defparam add_33937_7.INIT0 = 16'hf555;
    defparam add_33937_7.INIT1 = 16'hf555;
    defparam add_33937_7.INJECT1_0 = "NO";
    defparam add_33937_7.INJECT1_1 = "NO";
    CCU2D add_33937_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48771), .COUT(n48772));
    defparam add_33937_5.INIT0 = 16'hf555;
    defparam add_33937_5.INIT1 = 16'hf555;
    defparam add_33937_5.INJECT1_0 = "NO";
    defparam add_33937_5.INJECT1_1 = "NO";
    CCU2D add_33937_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48770), .COUT(n48771));
    defparam add_33937_3.INIT0 = 16'hf555;
    defparam add_33937_3.INIT1 = 16'hf555;
    defparam add_33937_3.INJECT1_0 = "NO";
    defparam add_33937_3.INJECT1_1 = "NO";
    CCU2D add_33937_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48770));
    defparam add_33937_1.INIT0 = 16'hF000;
    defparam add_33937_1.INIT1 = 16'ha666;
    defparam add_33937_1.INJECT1_0 = "NO";
    defparam add_33937_1.INJECT1_1 = "NO";
    PFUMX i37755 (.BLUT(n52955), .ALUT(n52956), .C0(bit_counter[1]), .Z(n52961));
    PFUMX i38965 (.BLUT(n54986), .ALUT(n54987), .C0(state[0]), .Z(state_2__N_104[1]));
    LUT4 i37751_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n52957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37751_3_lut.init = 16'hcaca;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47592), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47591), .COUT(n47592), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47590), .COUT(n47591), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47589), .COUT(n47590), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    PFUMX i38943 (.BLUT(n54952), .ALUT(n54953), .C0(state[1]), .Z(state_2__N_104[2]));
    PFUMX i38919 (.BLUT(n54916), .ALUT(n54917), .C0(state[1]), .Z(n52676));
    PFUMX i38917 (.BLUT(n54913), .ALUT(n54914), .C0(state[0]), .Z(n54915));
    PFUMX i38911 (.BLUT(n54904), .ALUT(n54905), .C0(state[1]), .Z(n54906));
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47588), .COUT(n47589), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U36 
//

module \WS2812(48000000,"111111111")_U36  (sclk_c, \port_status[12] , ws2813_out_c_12, 
            GND_net, \Q[12] , \RdAddress[12] );
    input sclk_c;
    output \port_status[12] ;
    output ws2813_out_c_12;
    input GND_net;
    input [23:0]\Q[12] ;
    output [8:0]\RdAddress[12] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_2220;
    wire [31:0]n9013;
    wire [31:0]n8837;
    
    wire n54706, n9012, n54596, sclk_c_enable_113, n54780, sclk_c_enable_114, 
        serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_118;
    wire [2:0]state_2__N_104;
    
    wire n47673;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n13696;
    wire [31:0]bit_counter_31__N_204;
    
    wire n47674, n53109, n53110, n53113, n47672, n53111, n53112, 
        n53114, n13731, n76, n8289, n103;
    wire [31:0]n447;
    
    wire n54944, n54943, n54649, n42582, n54650, n54587, n54712, 
        n69, n68;
    wire [6:0]n15073;
    
    wire sclk_c_enable_2038, n54794, n38412, sclk_c_enable_2005;
    wire [31:0]bit_counter_31__N_172;
    
    wire n54999, n54998, n35700, n53324, n53325, n53326, serial_N_437;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n35878;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_2069, n53101, n53102, n53103, n53104, n53105, 
        n53106, n53107, n53108;
    wire [8:0]n118;
    
    wire n53323, n53322, n53321, n53320, n52745, n35696, n53115, 
        n15, n14, n1, n1_adj_910, n54945, n55000, n47882, n47881, 
        n47880, n47879, n47878, n47877, n47876, n47875, n47874, 
        n47873, n47872, n47871, n47870, n47869, n47868, n47867, 
        n4, n47687, n47686, n47685, n47684, n47683, n47682, n48657, 
        n48656, n48655, n47817, n48654, n48653, n47816, n48652, 
        n48651, n48650, n48649, n48648, n48647, n48646, n48645, 
        n48644, n48643, n47815, n48642, n47681, n47680, n47814, 
        n47679, n47678, n48609, n48608, n48607, n48606, n48605, 
        n48604, n48603, n48602, n48601, n48600, n48599, n48598, 
        n48597, n48596, n48595, n48594, n47677, n47676, n47675;
    
    FD1P3AX delay_counter_i0_i0 (.D(n9013[0]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    LUT4 mux_2535_i9_4_lut (.A(n8837[8]), .B(n54706), .C(n9012), .D(n54596), 
         .Z(n9013[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i9_4_lut.init = 16'h303a;
    FD1P3AX status_77 (.D(n54780), .SP(sclk_c_enable_113), .CK(sclk_c), 
            .Q(\port_status[12] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_114), .CK(sclk_c), 
            .Q(ws2813_out_c_12)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_118), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_118), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_118), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_3126_5 (.A0(bit_counter[3]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47673), .COUT(n47674), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_5.INIT0 = 16'h5999;
    defparam add_3126_5.INIT1 = 16'h5999;
    defparam add_3126_5.INJECT1_0 = "NO";
    defparam add_3126_5.INJECT1_1 = "NO";
    L6MUX21 i37907 (.D0(n53109), .D1(n53110), .SD(bit_counter[2]), .Z(n53113));
    CCU2D add_3126_3 (.A0(bit_counter[1]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47672), .COUT(n47673), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_3.INIT0 = 16'h5999;
    defparam add_3126_3.INIT1 = 16'h5999;
    defparam add_3126_3.INJECT1_0 = "NO";
    defparam add_3126_3.INJECT1_1 = "NO";
    CCU2D add_3126_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13696), .C1(GND_net), .D1(GND_net), 
          .COUT(n47672), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_1.INIT0 = 16'hF000;
    defparam add_3126_1.INIT1 = 16'h5999;
    defparam add_3126_1.INJECT1_0 = "NO";
    defparam add_3126_1.INJECT1_1 = "NO";
    L6MUX21 i37908 (.D0(n53111), .D1(n53112), .SD(bit_counter[2]), .Z(n53114));
    LUT4 i38443_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .D(n13731), .Z(sclk_c_enable_118)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38443_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 mux_2535_i10_4_lut (.A(n76), .B(n54706), .C(n9012), .D(n54596), 
         .Z(n9013[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i10_4_lut.init = 16'h303a;
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13731), .Z(n8289)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 mux_2535_i13_4_lut (.A(n54596), .B(n54706), .C(n9012), .D(n103), 
         .Z(n9013[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i13_4_lut.init = 16'h3530;
    LUT4 mux_2525_i5_4_lut_4_lut_then_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13731), .Z(n54944)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2525_i5_4_lut_4_lut_then_4_lut.init = 16'he2e0;
    LUT4 mux_2525_i5_4_lut_4_lut_else_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13731), .Z(n54943)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2525_i5_4_lut_4_lut_else_4_lut.init = 16'hd0f0;
    LUT4 i1_2_lut_rep_646 (.A(state[2]), .B(n13731), .Z(n54649)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_646.init = 16'h4444;
    LUT4 i1_2_lut_rep_593_3_lut (.A(state[2]), .B(n13731), .C(state[1]), 
         .Z(n54596)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_593_3_lut.init = 16'h4040;
    LUT4 i38590_3_lut_rep_594_4_lut (.A(state[2]), .B(n13731), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2220)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38590_3_lut_rep_594_4_lut.init = 16'hfffb;
    LUT4 i37685_2_lut_rep_647 (.A(n42582), .B(n13696), .Z(n54650)) /* synthesis lut_function=(A (B)) */ ;
    defparam i37685_2_lut_rep_647.init = 16'h8888;
    LUT4 i1_2_lut_rep_584_3_lut (.A(n42582), .B(n13696), .C(state[1]), 
         .Z(n54587)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_584_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42582), .B(n13696), .C(n54712), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_709_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54712)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_709_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_584 (.A(state[2]), .B(state[1]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_584.init = 16'he0f0;
    LUT4 i1_2_lut_rep_703_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54706)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_703_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13731), 
         .Z(sclk_c_enable_114)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n15073[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_rep_680_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_2038)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_680_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_rep_791 (.A(state[2]), .B(state[0]), .Z(n54794)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_791.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_585 (.A(state[2]), .B(state[0]), .C(n13696), 
         .D(state[1]), .Z(n38412)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_585.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13696), 
         .D(state[1]), .Z(sclk_c_enable_2005)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_3_lut_adj_586 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_586.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_587 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_587.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_588 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_588.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_589 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_589.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_590 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_590.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_591 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_591.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_592 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_592.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_593 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_593.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_594 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_594.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_595 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_595.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_596 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_596.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_597 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_597.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_598 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_598.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_599 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_599.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_600 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_600.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_601 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_601.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_602 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_602.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_603 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_603.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_604 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_604.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_605 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_605.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_606 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_606.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_607 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_607.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_608 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_608.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_609 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_609.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_610 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_610.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_611 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_611.init = 16'h4040;
    LUT4 mux_2525_i3_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13731), .Z(n54999)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2525_i3_4_lut_then_4_lut.init = 16'hb1f0;
    LUT4 i1_2_lut_3_lut_adj_612 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_612.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_613 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_613.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_614 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_614.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_615 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_615.init = 16'h4040;
    LUT4 mux_2525_i3_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13696), .Z(n54998)) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2525_i3_4_lut_else_4_lut.init = 16'hb0f4;
    LUT4 i1_3_lut_4_lut (.A(n54587), .B(n54794), .C(n447[7]), .D(n54712), 
         .Z(n8837[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_616 (.A(n54587), .B(n54794), .C(n447[8]), 
         .D(n54712), .Z(n8837[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_616.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_617 (.A(n54587), .B(n54794), .C(n447[9]), 
         .D(n54712), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_617.init = 16'hf888;
    LUT4 i23508_4_lut (.A(sclk_c_enable_2220), .B(n54712), .C(n9012), 
         .D(n54596), .Z(n35700)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23508_4_lut.init = 16'haaa2;
    L6MUX21 i38120 (.D0(n53324), .D1(n53325), .SD(bit_counter[2]), .Z(n53326));
    FD1P3AX delay_counter_i0_i1 (.D(n9013[1]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n9013[3]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n9013[7]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n9013[8]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n9013[9]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n9013[12]), .SP(sclk_c_enable_2220), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i19520_1_lut_rep_777 (.A(state[2]), .Z(n54780)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i19520_1_lut_rep_777.init = 16'h5555;
    LUT4 i28939_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28939_3_lut_3_lut.init = 16'h5151;
    FD1P3IX pixel_i0 (.D(\Q[12] [0]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 mux_2395_i2_4_lut_4_lut (.A(n54706), .B(n54712), .C(n8289), .D(n13696), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2395_i2_4_lut_4_lut.init = 16'h5053;
    PFUMX i37903 (.BLUT(n53101), .ALUT(n53102), .C0(bit_counter[1]), .Z(n53109));
    PFUMX i37904 (.BLUT(n53103), .ALUT(n53104), .C0(bit_counter[1]), .Z(n53110));
    PFUMX i37905 (.BLUT(n53105), .ALUT(n53106), .C0(bit_counter[1]), .Z(n53111));
    PFUMX i37906 (.BLUT(n53107), .ALUT(n53108), .C0(bit_counter[1]), .Z(n53112));
    LUT4 i38400_2_lut_rep_838 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_2069)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38400_2_lut_rep_838.init = 16'h9999;
    LUT4 i23637_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35878)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23637_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_618 (.A(state[2]), .B(n42582), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_618.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_619 (.A(state[2]), .B(n42582), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_619.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_620 (.A(state[2]), .B(n42582), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_620.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_621 (.A(state[2]), .B(n42582), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_621.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_622 (.A(state[2]), .B(n42582), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_622.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_623 (.A(state[2]), .B(n42582), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_623.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_624 (.A(state[2]), .B(n42582), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_624.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_625 (.A(state[2]), .B(n42582), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_625.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_626 (.A(state[2]), .B(n42582), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_626.init = 16'h1010;
    LUT4 i38117_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38117_3_lut.init = 16'hcaca;
    LUT4 i38116_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38116_3_lut.init = 16'hcaca;
    LUT4 i38115_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38115_3_lut.init = 16'hcaca;
    LUT4 i38114_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38114_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54794), .B(state[1]), .C(n54650), .D(n54649), 
         .Z(n52745)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54650), .C(n13731), .D(n54794), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    LUT4 i23484_2_lut_4_lut (.A(n54649), .B(state[0]), .C(state[1]), .D(n9012), 
         .Z(n35696)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23484_2_lut_4_lut.init = 16'hfd00;
    LUT4 i37902_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37902_3_lut.init = 16'hcaca;
    LUT4 i37901_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37901_3_lut.init = 16'hcaca;
    LUT4 i37900_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37900_3_lut.init = 16'hcaca;
    LUT4 i37899_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37899_3_lut.init = 16'hcaca;
    LUT4 i37898_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37898_3_lut.init = 16'hcaca;
    LUT4 i37897_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37897_3_lut.init = 16'hcaca;
    LUT4 i37896_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37896_3_lut.init = 16'hcaca;
    LUT4 i37895_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37895_3_lut.init = 16'hcaca;
    L6MUX21 i37909 (.D0(n53113), .D1(n53114), .SD(bit_counter[3]), .Z(n53115));
    PFUMX i38118 (.BLUT(n53320), .ALUT(n53321), .C0(bit_counter[1]), .Z(n53324));
    PFUMX i38119 (.BLUT(n53322), .ALUT(n53323), .C0(bit_counter[1]), .Z(n53325));
    LUT4 mux_2535_i1_4_lut (.A(n69), .B(n15073[0]), .C(n9012), .D(n52745), 
         .Z(n9013[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i1_4_lut.init = 16'hcfca;
    LUT4 i2547_3_lut (.A(state[2]), .B(state[1]), .C(n13731), .Z(n9012)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2547_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[2]), .C(n14), .D(cur_pixel[8]), 
         .Z(n42582)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[3]), .B(cur_pixel[5]), .C(cur_pixel[7]), 
         .D(cur_pixel[4]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[6]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    FD1P3IX pixel_i23 (.D(\Q[12] [23]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[12] [22]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[12] [21]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[12] [20]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[12] [19]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[12] [18]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[12] [17]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[12] [16]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[12] [15]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[12] [14]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[12] [13]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[12] [12]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[12] [11]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[12] [10]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[12] [9]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[12] [8]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[12] [7]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[12] [6]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[12] [5]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[12] [4]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[12] [3]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[12] [2]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[12] [1]), .SP(sclk_c_enable_2038), .CD(n35878), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2005), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2038), 
            .CD(n35878), .CK(sclk_c), .Q(\RdAddress[12] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53115), .B(n53326), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_2069), .CD(n35878), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_910), .SP(sclk_c_enable_2069), .CD(n35878), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_2069), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 mux_2395_i1_4_lut (.A(n54650), .B(n54706), .C(n8289), .D(n54712), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2395_i1_4_lut.init = 16'h3f3a;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2220), 
            .CD(n35700), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2220), .CD(n35700), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2220), .CD(n35700), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54945), .SP(sclk_c_enable_2220), .CD(n35696), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n55000), .SP(sclk_c_enable_2220), .CD(n35696), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=267, LSE_RLINE=267 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47882), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47881), .COUT(n47882), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47880), .COUT(n47881), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47879), .COUT(n47880), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47878), .COUT(n47879), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47877), .COUT(n47878), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47876), .COUT(n47877), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47875), .COUT(n47876), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47874), .COUT(n47875), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47873), .COUT(n47874), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    LUT4 i28780_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28780_2_lut.init = 16'hbbbb;
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47872), .COUT(n47873), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47871), .COUT(n47872), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47870), .COUT(n47871), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47869), .COUT(n47870), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i28779_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_910)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28779_2_lut.init = 16'hbbbb;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47868), .COUT(n47869), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47867), .COUT(n47868), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47867), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 mux_2535_i2_4_lut (.A(n68), .B(n15073[0]), .C(n9012), .D(n52745), 
         .Z(n9013[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2535_i4_4_lut (.A(n38412), .B(n54706), .C(n9012), .D(n4), 
         .Z(n9013[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42582), .B(n54596), .C(n447[3]), .D(n54712), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2535_i8_4_lut (.A(n8837[7]), .B(n54706), .C(n9012), .D(n54596), 
         .Z(n9013[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2535_i8_4_lut.init = 16'h303a;
    PFUMX i38973 (.BLUT(n54998), .ALUT(n54999), .C0(state[1]), .Z(n55000));
    CCU2D add_3126_33 (.A0(bit_counter[31]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47687), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_33.INIT0 = 16'h5999;
    defparam add_3126_33.INIT1 = 16'h0000;
    defparam add_3126_33.INJECT1_0 = "NO";
    defparam add_3126_33.INJECT1_1 = "NO";
    CCU2D add_3126_31 (.A0(bit_counter[29]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47686), .COUT(n47687), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_31.INIT0 = 16'h5999;
    defparam add_3126_31.INIT1 = 16'h5999;
    defparam add_3126_31.INJECT1_0 = "NO";
    defparam add_3126_31.INJECT1_1 = "NO";
    CCU2D add_3126_29 (.A0(bit_counter[27]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47685), .COUT(n47686), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_29.INIT0 = 16'h5999;
    defparam add_3126_29.INIT1 = 16'h5999;
    defparam add_3126_29.INJECT1_0 = "NO";
    defparam add_3126_29.INJECT1_1 = "NO";
    CCU2D add_3126_27 (.A0(bit_counter[25]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47684), .COUT(n47685), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_27.INIT0 = 16'h5999;
    defparam add_3126_27.INIT1 = 16'h5999;
    defparam add_3126_27.INJECT1_0 = "NO";
    defparam add_3126_27.INJECT1_1 = "NO";
    CCU2D add_3126_25 (.A0(bit_counter[23]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47683), .COUT(n47684), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_25.INIT0 = 16'h5999;
    defparam add_3126_25.INIT1 = 16'h5999;
    defparam add_3126_25.INJECT1_0 = "NO";
    defparam add_3126_25.INJECT1_1 = "NO";
    CCU2D add_3126_23 (.A0(bit_counter[21]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47682), .COUT(n47683), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_23.INIT0 = 16'h5999;
    defparam add_3126_23.INIT1 = 16'h5999;
    defparam add_3126_23.INJECT1_0 = "NO";
    defparam add_3126_23.INJECT1_1 = "NO";
    CCU2D add_33908_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48657), 
          .S0(n13731));
    defparam add_33908_cout.INIT0 = 16'h0000;
    defparam add_33908_cout.INIT1 = 16'h0000;
    defparam add_33908_cout.INJECT1_0 = "NO";
    defparam add_33908_cout.INJECT1_1 = "NO";
    CCU2D add_33908_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48656), .COUT(n48657));
    defparam add_33908_31.INIT0 = 16'hf555;
    defparam add_33908_31.INIT1 = 16'h5555;
    defparam add_33908_31.INJECT1_0 = "NO";
    defparam add_33908_31.INJECT1_1 = "NO";
    CCU2D add_33908_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48655), .COUT(n48656));
    defparam add_33908_29.INIT0 = 16'hf555;
    defparam add_33908_29.INIT1 = 16'hf555;
    defparam add_33908_29.INJECT1_0 = "NO";
    defparam add_33908_29.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47817), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_33908_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48654), .COUT(n48655));
    defparam add_33908_27.INIT0 = 16'hf555;
    defparam add_33908_27.INIT1 = 16'hf555;
    defparam add_33908_27.INJECT1_0 = "NO";
    defparam add_33908_27.INJECT1_1 = "NO";
    CCU2D add_33908_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48653), .COUT(n48654));
    defparam add_33908_25.INIT0 = 16'hf555;
    defparam add_33908_25.INIT1 = 16'hf555;
    defparam add_33908_25.INJECT1_0 = "NO";
    defparam add_33908_25.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47816), .COUT(n47817), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_33908_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48652), .COUT(n48653));
    defparam add_33908_23.INIT0 = 16'hf555;
    defparam add_33908_23.INIT1 = 16'hf555;
    defparam add_33908_23.INJECT1_0 = "NO";
    defparam add_33908_23.INJECT1_1 = "NO";
    CCU2D add_33908_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48651), .COUT(n48652));
    defparam add_33908_21.INIT0 = 16'hf555;
    defparam add_33908_21.INIT1 = 16'hf555;
    defparam add_33908_21.INJECT1_0 = "NO";
    defparam add_33908_21.INJECT1_1 = "NO";
    CCU2D add_33908_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48650), .COUT(n48651));
    defparam add_33908_19.INIT0 = 16'hf555;
    defparam add_33908_19.INIT1 = 16'hf555;
    defparam add_33908_19.INJECT1_0 = "NO";
    defparam add_33908_19.INJECT1_1 = "NO";
    CCU2D add_33908_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48649), .COUT(n48650));
    defparam add_33908_17.INIT0 = 16'hf555;
    defparam add_33908_17.INIT1 = 16'hf555;
    defparam add_33908_17.INJECT1_0 = "NO";
    defparam add_33908_17.INJECT1_1 = "NO";
    CCU2D add_33908_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48648), .COUT(n48649));
    defparam add_33908_15.INIT0 = 16'hf555;
    defparam add_33908_15.INIT1 = 16'hf555;
    defparam add_33908_15.INJECT1_0 = "NO";
    defparam add_33908_15.INJECT1_1 = "NO";
    CCU2D add_33908_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48647), .COUT(n48648));
    defparam add_33908_13.INIT0 = 16'hf555;
    defparam add_33908_13.INIT1 = 16'hf555;
    defparam add_33908_13.INJECT1_0 = "NO";
    defparam add_33908_13.INJECT1_1 = "NO";
    CCU2D add_33908_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48646), .COUT(n48647));
    defparam add_33908_11.INIT0 = 16'hf555;
    defparam add_33908_11.INIT1 = 16'hf555;
    defparam add_33908_11.INJECT1_0 = "NO";
    defparam add_33908_11.INJECT1_1 = "NO";
    CCU2D add_33908_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48645), .COUT(n48646));
    defparam add_33908_9.INIT0 = 16'hf555;
    defparam add_33908_9.INIT1 = 16'hf555;
    defparam add_33908_9.INJECT1_0 = "NO";
    defparam add_33908_9.INJECT1_1 = "NO";
    CCU2D add_33908_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48644), .COUT(n48645));
    defparam add_33908_7.INIT0 = 16'hf555;
    defparam add_33908_7.INIT1 = 16'hf555;
    defparam add_33908_7.INJECT1_0 = "NO";
    defparam add_33908_7.INJECT1_1 = "NO";
    CCU2D add_33908_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48643), .COUT(n48644));
    defparam add_33908_5.INIT0 = 16'hf555;
    defparam add_33908_5.INIT1 = 16'hf555;
    defparam add_33908_5.INJECT1_0 = "NO";
    defparam add_33908_5.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47815), .COUT(n47816), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_33908_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48642), .COUT(n48643));
    defparam add_33908_3.INIT0 = 16'hf555;
    defparam add_33908_3.INIT1 = 16'hf555;
    defparam add_33908_3.INJECT1_0 = "NO";
    defparam add_33908_3.INJECT1_1 = "NO";
    CCU2D add_3126_21 (.A0(bit_counter[19]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47681), .COUT(n47682), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_21.INIT0 = 16'h5999;
    defparam add_3126_21.INIT1 = 16'h5999;
    defparam add_3126_21.INJECT1_0 = "NO";
    defparam add_3126_21.INJECT1_1 = "NO";
    CCU2D add_33908_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48642));
    defparam add_33908_1.INIT0 = 16'hF000;
    defparam add_33908_1.INIT1 = 16'ha666;
    defparam add_33908_1.INJECT1_0 = "NO";
    defparam add_33908_1.INJECT1_1 = "NO";
    CCU2D add_3126_19 (.A0(bit_counter[17]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47680), .COUT(n47681), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_19.INIT0 = 16'h5999;
    defparam add_3126_19.INIT1 = 16'h5999;
    defparam add_3126_19.INJECT1_0 = "NO";
    defparam add_3126_19.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47814), .COUT(n47815), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    PFUMX i38937 (.BLUT(n54943), .ALUT(n54944), .C0(state[0]), .Z(n54945));
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47814), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3126_17 (.A0(bit_counter[15]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47679), .COUT(n47680), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_17.INIT0 = 16'h5999;
    defparam add_3126_17.INIT1 = 16'h5999;
    defparam add_3126_17.INJECT1_0 = "NO";
    defparam add_3126_17.INJECT1_1 = "NO";
    CCU2D add_3126_15 (.A0(bit_counter[13]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47678), .COUT(n47679), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_15.INIT0 = 16'h5999;
    defparam add_3126_15.INIT1 = 16'h5999;
    defparam add_3126_15.INJECT1_0 = "NO";
    defparam add_3126_15.INJECT1_1 = "NO";
    CCU2D add_33909_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48609), 
          .S0(n13696));
    defparam add_33909_cout.INIT0 = 16'h0000;
    defparam add_33909_cout.INIT1 = 16'h0000;
    defparam add_33909_cout.INJECT1_0 = "NO";
    defparam add_33909_cout.INJECT1_1 = "NO";
    CCU2D add_33909_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48608), .COUT(n48609));
    defparam add_33909_31.INIT0 = 16'hf555;
    defparam add_33909_31.INIT1 = 16'h5555;
    defparam add_33909_31.INJECT1_0 = "NO";
    defparam add_33909_31.INJECT1_1 = "NO";
    CCU2D add_33909_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48607), .COUT(n48608));
    defparam add_33909_29.INIT0 = 16'hf555;
    defparam add_33909_29.INIT1 = 16'hf555;
    defparam add_33909_29.INJECT1_0 = "NO";
    defparam add_33909_29.INJECT1_1 = "NO";
    CCU2D add_33909_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48606), .COUT(n48607));
    defparam add_33909_27.INIT0 = 16'hf555;
    defparam add_33909_27.INIT1 = 16'hf555;
    defparam add_33909_27.INJECT1_0 = "NO";
    defparam add_33909_27.INJECT1_1 = "NO";
    CCU2D add_33909_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48605), .COUT(n48606));
    defparam add_33909_25.INIT0 = 16'hf555;
    defparam add_33909_25.INIT1 = 16'hf555;
    defparam add_33909_25.INJECT1_0 = "NO";
    defparam add_33909_25.INJECT1_1 = "NO";
    CCU2D add_33909_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48604), .COUT(n48605));
    defparam add_33909_23.INIT0 = 16'hf555;
    defparam add_33909_23.INIT1 = 16'hf555;
    defparam add_33909_23.INJECT1_0 = "NO";
    defparam add_33909_23.INJECT1_1 = "NO";
    CCU2D add_33909_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48603), .COUT(n48604));
    defparam add_33909_21.INIT0 = 16'hf555;
    defparam add_33909_21.INIT1 = 16'hf555;
    defparam add_33909_21.INJECT1_0 = "NO";
    defparam add_33909_21.INJECT1_1 = "NO";
    CCU2D add_33909_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48602), .COUT(n48603));
    defparam add_33909_19.INIT0 = 16'hf555;
    defparam add_33909_19.INIT1 = 16'hf555;
    defparam add_33909_19.INJECT1_0 = "NO";
    defparam add_33909_19.INJECT1_1 = "NO";
    CCU2D add_33909_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48601), .COUT(n48602));
    defparam add_33909_17.INIT0 = 16'hf555;
    defparam add_33909_17.INIT1 = 16'hf555;
    defparam add_33909_17.INJECT1_0 = "NO";
    defparam add_33909_17.INJECT1_1 = "NO";
    CCU2D add_33909_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48600), .COUT(n48601));
    defparam add_33909_15.INIT0 = 16'hf555;
    defparam add_33909_15.INIT1 = 16'hf555;
    defparam add_33909_15.INJECT1_0 = "NO";
    defparam add_33909_15.INJECT1_1 = "NO";
    CCU2D add_33909_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48599), .COUT(n48600));
    defparam add_33909_13.INIT0 = 16'hf555;
    defparam add_33909_13.INIT1 = 16'hf555;
    defparam add_33909_13.INJECT1_0 = "NO";
    defparam add_33909_13.INJECT1_1 = "NO";
    CCU2D add_33909_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48598), .COUT(n48599));
    defparam add_33909_11.INIT0 = 16'hf555;
    defparam add_33909_11.INIT1 = 16'hf555;
    defparam add_33909_11.INJECT1_0 = "NO";
    defparam add_33909_11.INJECT1_1 = "NO";
    CCU2D add_33909_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48597), .COUT(n48598));
    defparam add_33909_9.INIT0 = 16'hf555;
    defparam add_33909_9.INIT1 = 16'hf555;
    defparam add_33909_9.INJECT1_0 = "NO";
    defparam add_33909_9.INJECT1_1 = "NO";
    CCU2D add_33909_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48596), .COUT(n48597));
    defparam add_33909_7.INIT0 = 16'hf555;
    defparam add_33909_7.INIT1 = 16'hf555;
    defparam add_33909_7.INJECT1_0 = "NO";
    defparam add_33909_7.INJECT1_1 = "NO";
    CCU2D add_33909_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48595), .COUT(n48596));
    defparam add_33909_5.INIT0 = 16'hf555;
    defparam add_33909_5.INIT1 = 16'hf555;
    defparam add_33909_5.INJECT1_0 = "NO";
    defparam add_33909_5.INJECT1_1 = "NO";
    CCU2D add_33909_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48594), .COUT(n48595));
    defparam add_33909_3.INIT0 = 16'hf555;
    defparam add_33909_3.INIT1 = 16'hf555;
    defparam add_33909_3.INJECT1_0 = "NO";
    defparam add_33909_3.INJECT1_1 = "NO";
    CCU2D add_3126_13 (.A0(bit_counter[11]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47677), .COUT(n47678), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_13.INIT0 = 16'h5999;
    defparam add_3126_13.INIT1 = 16'h5999;
    defparam add_3126_13.INJECT1_0 = "NO";
    defparam add_3126_13.INJECT1_1 = "NO";
    CCU2D add_33909_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48594));
    defparam add_33909_1.INIT0 = 16'hF000;
    defparam add_33909_1.INIT1 = 16'ha666;
    defparam add_33909_1.INJECT1_0 = "NO";
    defparam add_33909_1.INJECT1_1 = "NO";
    CCU2D add_3126_11 (.A0(bit_counter[9]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47676), .COUT(n47677), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_11.INIT0 = 16'h5999;
    defparam add_3126_11.INIT1 = 16'h5999;
    defparam add_3126_11.INJECT1_0 = "NO";
    defparam add_3126_11.INJECT1_1 = "NO";
    CCU2D add_3126_9 (.A0(bit_counter[7]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47675), .COUT(n47676), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_9.INIT0 = 16'h5999;
    defparam add_3126_9.INIT1 = 16'h5999;
    defparam add_3126_9.INJECT1_0 = "NO";
    defparam add_3126_9.INJECT1_1 = "NO";
    CCU2D add_3126_7 (.A0(bit_counter[5]), .B0(n13696), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13696), .C1(GND_net), 
          .D1(GND_net), .CIN(n47674), .COUT(n47675), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3126_7.INIT0 = 16'h5999;
    defparam add_3126_7.INIT1 = 16'h5999;
    defparam add_3126_7.INJECT1_0 = "NO";
    defparam add_3126_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U23 
//

module \WS2812(48000000,"111111111")_U23  (sclk_c, \port_status[5] , ws2813_out_c_5, 
            GND_net, \Q[5] , \RdAddress[5] );
    input sclk_c;
    output \port_status[5] ;
    output ws2813_out_c_5;
    input GND_net;
    input [23:0]\Q[5] ;
    output [8:0]\RdAddress[5] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_921;
    wire [31:0]n6832;
    
    wire sclk_c_enable_52, n54817, sclk_c_enable_53, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_57;
    wire [2:0]state_2__N_104;
    
    wire n47671;
    wire [31:0]n447;
    
    wire n47670, n13241, n9936;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1202, n35213, n54923, n13206, n54922;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1188;
    wire [8:0]cur_pixel_8__N_107;
    
    wire n54981, n54980, n53275, n53276;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53277, sclk_c_enable_1203;
    wire [31:0]bit_counter_31__N_172;
    
    wire n1, n1_adj_909, n35035, n35031, n54982, n54924, n48561, 
        n47669, n48560, n54670, n54556, n48559, n54607, n54825, 
        n54684;
    wire [31:0]n6656;
    
    wire n76, serial_N_437, n48558, n69, n68;
    wire [6:0]n15006;
    
    wire n54724, n39343;
    wire [31:0]bit_counter_31__N_204;
    
    wire n52996, n52997, n53004, n52998, n52999, n53005, n53000, 
        n53001, n53006, n53002, n53003, n53007, n48557, n47668, 
        n48556, n47667, n42588;
    wire [8:0]n118;
    
    wire n48555, n48554, n48553, n47666, n47665, n48552, n47664, 
        n47663, n48551, n48550, n15, n14, n48549, n48548, n48547, 
        n48546, n47662, n47661, n6831, n53010, n54619, n53274, 
        n53273, n47660, n53272, n53271, n47659, n47658, n47657, 
        n47656, n47654, n47653, n47652, n47651, n52733, n53008, 
        n53009, n48162, n48161, n48160, n48159, n48158, n48157, 
        n48156, n48155, n48154, n48153, n48152, n48151, n48150, 
        n48149, n48148, n48147, n4, n103, n48338, n48337, n48336, 
        n48335, n48334, n48333, n48332, n48331, n48330, n48329, 
        n48328, n48327, n48326, n48325, n48324, n48323;
    
    FD1P3AX delay_counter_i0_i0 (.D(n6832[0]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54817), .SP(sclk_c_enable_52), .CK(sclk_c), 
            .Q(\port_status[5] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_53), .CK(sclk_c), 
            .Q(ws2813_out_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_57), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_57), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_57), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47671), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47670), .COUT(n47671), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    LUT4 i38447_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13241), .Z(sclk_c_enable_57)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38447_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13241), .Z(n9936)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    FD1P3IX pixel_i23 (.D(\Q[5] [23]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[5] [22]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[5] [21]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[5] [20]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[5] [19]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[5] [18]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[5] [17]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[5] [16]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[5] [15]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[5] [14]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[5] [13]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[5] [12]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[5] [11]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[5] [10]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[5] [9]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[5] [8]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[5] [7]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[5] [6]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[5] [5]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[5] [4]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    LUT4 mux_2042_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13241), .Z(n54923)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2042_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2042_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13206), .Z(n54922)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2042_i3_4_lut_else_4_lut.init = 16'hd0f2;
    FD1P3IX pixel_i3 (.D(\Q[5] [3]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[5] [2]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[5] [1]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    LUT4 mux_2042_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13241), .Z(n54981)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2042_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2042_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13241), .Z(n54980)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2042_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    L6MUX21 i38071 (.D0(n53275), .D1(n53276), .SD(bit_counter[2]), .Z(n53277));
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1203), .CD(n35213), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_909), .SP(sclk_c_enable_1203), .CD(n35213), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_921), 
            .CD(n35035), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_921), .CD(n35035), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_921), .CD(n35035), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54982), .SP(sclk_c_enable_921), .CD(n35031), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54924), .SP(sclk_c_enable_921), .CD(n35031), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    CCU2D add_33912_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48561), 
          .S0(n13241));
    defparam add_33912_cout.INIT0 = 16'h0000;
    defparam add_33912_cout.INIT1 = 16'h0000;
    defparam add_33912_cout.INJECT1_0 = "NO";
    defparam add_33912_cout.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47669), .COUT(n47670), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_33912_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48560), .COUT(n48561));
    defparam add_33912_31.INIT0 = 16'hf555;
    defparam add_33912_31.INIT1 = 16'h5555;
    defparam add_33912_31.INJECT1_0 = "NO";
    defparam add_33912_31.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_667 (.A(state[2]), .B(n13241), .Z(n54670)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_667.init = 16'h4444;
    LUT4 i1_2_lut_rep_553_3_lut (.A(state[2]), .B(n13241), .C(state[1]), 
         .Z(n54556)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_553_3_lut.init = 16'h4040;
    LUT4 i38613_3_lut_rep_557_4_lut (.A(state[2]), .B(n13241), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_921)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38613_3_lut_rep_557_4_lut.init = 16'hfffb;
    FD1P3AX delay_counter_i0_i1 (.D(n6832[1]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n6832[3]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n6832[7]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n6832[8]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n6832[9]), .SP(sclk_c_enable_921), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n6832[12]), .SP(sclk_c_enable_921), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    CCU2D add_33912_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48559), .COUT(n48560));
    defparam add_33912_29.INIT0 = 16'hf555;
    defparam add_33912_29.INIT1 = 16'hf555;
    defparam add_33912_29.INJECT1_0 = "NO";
    defparam add_33912_29.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(n54607), .B(n54825), .C(n447[7]), .D(n54684), 
         .Z(n6656[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_541 (.A(n54607), .B(n54825), .C(n447[8]), 
         .D(n54684), .Z(n6656[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_541.init = 16'hf888;
    LUT4 i38430_2_lut_rep_812 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1203)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38430_2_lut_rep_812.init = 16'h9999;
    LUT4 i1_3_lut_4_lut_adj_542 (.A(n54607), .B(n54825), .C(n447[9]), 
         .D(n54684), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_542.init = 16'hf888;
    LUT4 i27151_1_lut_rep_814 (.A(state[2]), .Z(n54817)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27151_1_lut_rep_814.init = 16'h5555;
    LUT4 i28902_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28902_3_lut_3_lut.init = 16'h5151;
    CCU2D add_33912_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48558), .COUT(n48559));
    defparam add_33912_27.INIT0 = 16'hf555;
    defparam add_33912_27.INIT1 = 16'hf555;
    defparam add_33912_27.INJECT1_0 = "NO";
    defparam add_33912_27.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_681_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54684)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_681_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_543 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_543.init = 16'he0f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13241), 
         .Z(sclk_c_enable_53)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i23064_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35213)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23064_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_724_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1202)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_724_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n15006[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_721_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54724)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_721_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_822 (.A(state[0]), .B(state[2]), .Z(n54825)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_822.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_544 (.A(state[0]), .B(state[2]), .C(n13206), 
         .D(state[1]), .Z(n39343)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_544.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13206), 
         .D(state[1]), .Z(sclk_c_enable_1188)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_545 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_545.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_546 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_546.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_547 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_547.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_548 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_548.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_549 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_549.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_550 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_550.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_551 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_551.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_552 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_552.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_553 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_553.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_554 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_554.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_555 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_555.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_556 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_556.init = 16'h2020;
    PFUMX i37798 (.BLUT(n52996), .ALUT(n52997), .C0(bit_counter[1]), .Z(n53004));
    LUT4 i1_2_lut_3_lut_adj_557 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_557.init = 16'h2020;
    PFUMX i37799 (.BLUT(n52998), .ALUT(n52999), .C0(bit_counter[1]), .Z(n53005));
    LUT4 i1_2_lut_3_lut_adj_558 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_558.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_559 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_559.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_560 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_560.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_561 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_561.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_562 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_562.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_563 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_563.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_564 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_564.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_565 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_565.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_566 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_566.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_567 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_567.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_568 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_568.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_569 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_569.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_570 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_570.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_571 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_571.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_572 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_572.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_573 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_573.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_574 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_574.init = 16'h2020;
    PFUMX i37800 (.BLUT(n53000), .ALUT(n53001), .C0(bit_counter[1]), .Z(n53006));
    PFUMX i37801 (.BLUT(n53002), .ALUT(n53003), .C0(bit_counter[1]), .Z(n53007));
    FD1P3IX pixel_i0 (.D(\Q[5] [0]), .SP(sclk_c_enable_1202), .CD(n35213), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1188), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1202), 
            .CD(n35213), .CK(sclk_c), .Q(\RdAddress[5] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1203), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=190, LSE_RLINE=190 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 mux_2764_i2_4_lut_4_lut (.A(n54724), .B(n54684), .C(n9936), .D(n13206), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2764_i2_4_lut_4_lut.init = 16'h5053;
    CCU2D add_33912_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48557), .COUT(n48558));
    defparam add_33912_25.INIT0 = 16'hf555;
    defparam add_33912_25.INIT1 = 16'hf555;
    defparam add_33912_25.INJECT1_0 = "NO";
    defparam add_33912_25.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47668), .COUT(n47669), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_33912_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48556), .COUT(n48557));
    defparam add_33912_23.INIT0 = 16'hf555;
    defparam add_33912_23.INIT1 = 16'hf555;
    defparam add_33912_23.INJECT1_0 = "NO";
    defparam add_33912_23.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47667), .COUT(n47668), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_575 (.A(state[2]), .B(n42588), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_575.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_576 (.A(state[2]), .B(n42588), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_576.init = 16'h1010;
    CCU2D add_33912_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48555), .COUT(n48556));
    defparam add_33912_21.INIT0 = 16'hf555;
    defparam add_33912_21.INIT1 = 16'hf555;
    defparam add_33912_21.INJECT1_0 = "NO";
    defparam add_33912_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_577 (.A(state[2]), .B(n42588), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_577.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_578 (.A(state[2]), .B(n42588), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_578.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_579 (.A(state[2]), .B(n42588), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_579.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_580 (.A(state[2]), .B(n42588), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_580.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_581 (.A(state[2]), .B(n42588), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_581.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_582 (.A(state[2]), .B(n42588), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_582.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_583 (.A(state[2]), .B(n42588), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_583.init = 16'h1010;
    CCU2D add_33912_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48554), .COUT(n48555));
    defparam add_33912_19.INIT0 = 16'hf555;
    defparam add_33912_19.INIT1 = 16'hf555;
    defparam add_33912_19.INJECT1_0 = "NO";
    defparam add_33912_19.INJECT1_1 = "NO";
    CCU2D add_33912_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48553), .COUT(n48554));
    defparam add_33912_17.INIT0 = 16'hf555;
    defparam add_33912_17.INIT1 = 16'hf555;
    defparam add_33912_17.INJECT1_0 = "NO";
    defparam add_33912_17.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47666), .COUT(n47667), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47665), .COUT(n47666), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_33912_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48552), .COUT(n48553));
    defparam add_33912_15.INIT0 = 16'hf555;
    defparam add_33912_15.INIT1 = 16'hf555;
    defparam add_33912_15.INJECT1_0 = "NO";
    defparam add_33912_15.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47664), .COUT(n47665), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47663), .COUT(n47664), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_33912_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48551), .COUT(n48552));
    defparam add_33912_13.INIT0 = 16'hf555;
    defparam add_33912_13.INIT1 = 16'hf555;
    defparam add_33912_13.INJECT1_0 = "NO";
    defparam add_33912_13.INJECT1_1 = "NO";
    CCU2D add_33912_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48550), .COUT(n48551));
    defparam add_33912_11.INIT0 = 16'hf555;
    defparam add_33912_11.INIT1 = 16'hf555;
    defparam add_33912_11.INJECT1_0 = "NO";
    defparam add_33912_11.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[2]), .C(n14), .D(cur_pixel[8]), 
         .Z(n42588)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[3]), .B(cur_pixel[5]), .C(cur_pixel[7]), 
         .D(cur_pixel[4]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    CCU2D add_33912_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48549), .COUT(n48550));
    defparam add_33912_9.INIT0 = 16'hf555;
    defparam add_33912_9.INIT1 = 16'hf555;
    defparam add_33912_9.INJECT1_0 = "NO";
    defparam add_33912_9.INJECT1_1 = "NO";
    CCU2D add_33912_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48548), .COUT(n48549));
    defparam add_33912_7.INIT0 = 16'hf555;
    defparam add_33912_7.INIT1 = 16'hf555;
    defparam add_33912_7.INJECT1_0 = "NO";
    defparam add_33912_7.INJECT1_1 = "NO";
    LUT4 i5_3_lut (.A(cur_pixel[6]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    CCU2D add_33912_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48547), .COUT(n48548));
    defparam add_33912_5.INIT0 = 16'hf555;
    defparam add_33912_5.INIT1 = 16'hf555;
    defparam add_33912_5.INJECT1_0 = "NO";
    defparam add_33912_5.INJECT1_1 = "NO";
    CCU2D add_33912_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48546), .COUT(n48547));
    defparam add_33912_3.INIT0 = 16'hf555;
    defparam add_33912_3.INIT1 = 16'hf555;
    defparam add_33912_3.INJECT1_0 = "NO";
    defparam add_33912_3.INJECT1_1 = "NO";
    CCU2D add_33912_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48546));
    defparam add_33912_1.INIT0 = 16'hF000;
    defparam add_33912_1.INIT1 = 16'ha666;
    defparam add_33912_1.INJECT1_0 = "NO";
    defparam add_33912_1.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47662), .COUT(n47663), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47661), .COUT(n47662), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    LUT4 i22819_2_lut_4_lut (.A(n54670), .B(state[0]), .C(state[1]), .D(n6831), 
         .Z(n35031)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i22819_2_lut_4_lut.init = 16'hfd00;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53010), .B(n53277), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2764_i1_4_lut (.A(n54619), .B(n54724), .C(n9936), .D(n54684), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2764_i1_4_lut.init = 16'h3f3a;
    LUT4 i2064_3_lut (.A(state[2]), .B(state[1]), .C(n13241), .Z(n6831)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2064_3_lut.init = 16'ha8a8;
    LUT4 i38068_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38068_3_lut.init = 16'hcaca;
    LUT4 i38067_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38067_3_lut.init = 16'hcaca;
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47660), .COUT(n47661), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    LUT4 i38066_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38066_3_lut.init = 16'hcaca;
    LUT4 i38065_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38065_3_lut.init = 16'hcaca;
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47659), .COUT(n47660), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i28645_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28645_2_lut.init = 16'hbbbb;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47658), .COUT(n47659), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i28673_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_909)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28673_2_lut.init = 16'hbbbb;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47657), .COUT(n47658), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47656), .COUT(n47657), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47656), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47654), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47653), .COUT(n47654), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47652), .COUT(n47653), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47651), .COUT(n47652), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47651), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54825), .B(state[1]), .C(n54619), .D(n54670), 
         .Z(n52733)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    L6MUX21 i37804 (.D0(n53008), .D1(n53009), .SD(bit_counter[3]), .Z(n53010));
    LUT4 i22843_4_lut (.A(sclk_c_enable_921), .B(n54684), .C(n6831), .D(n54556), 
         .Z(n35035)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22843_4_lut.init = 16'haaa2;
    PFUMX i38069 (.BLUT(n53271), .ALUT(n53272), .C0(bit_counter[1]), .Z(n53275));
    PFUMX i38070 (.BLUT(n53273), .ALUT(n53274), .C0(bit_counter[1]), .Z(n53276));
    L6MUX21 i37802 (.D0(n53004), .D1(n53005), .SD(bit_counter[2]), .Z(n53008));
    L6MUX21 i37803 (.D0(n53006), .D1(n53007), .SD(bit_counter[2]), .Z(n53009));
    LUT4 i37797_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37797_3_lut.init = 16'hcaca;
    LUT4 i37796_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37796_3_lut.init = 16'hcaca;
    LUT4 i37795_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37795_3_lut.init = 16'hcaca;
    LUT4 i37794_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37794_3_lut.init = 16'hcaca;
    LUT4 i37793_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37793_3_lut.init = 16'hcaca;
    LUT4 i37792_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37792_3_lut.init = 16'hcaca;
    LUT4 i37791_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37791_3_lut.init = 16'hcaca;
    LUT4 i37790_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37790_3_lut.init = 16'hcaca;
    LUT4 mux_2052_i1_4_lut (.A(n69), .B(n15006[0]), .C(n6831), .D(n52733), 
         .Z(n6832[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i1_4_lut.init = 16'hcfca;
    CCU2D add_33919_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48162), 
          .S0(n13206));
    defparam add_33919_cout.INIT0 = 16'h0000;
    defparam add_33919_cout.INIT1 = 16'h0000;
    defparam add_33919_cout.INJECT1_0 = "NO";
    defparam add_33919_cout.INJECT1_1 = "NO";
    CCU2D add_33919_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48161), .COUT(n48162));
    defparam add_33919_31.INIT0 = 16'hf555;
    defparam add_33919_31.INIT1 = 16'h5555;
    defparam add_33919_31.INJECT1_0 = "NO";
    defparam add_33919_31.INJECT1_1 = "NO";
    CCU2D add_33919_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48160), .COUT(n48161));
    defparam add_33919_29.INIT0 = 16'hf555;
    defparam add_33919_29.INIT1 = 16'hf555;
    defparam add_33919_29.INJECT1_0 = "NO";
    defparam add_33919_29.INJECT1_1 = "NO";
    CCU2D add_33919_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48159), .COUT(n48160));
    defparam add_33919_27.INIT0 = 16'hf555;
    defparam add_33919_27.INIT1 = 16'hf555;
    defparam add_33919_27.INJECT1_0 = "NO";
    defparam add_33919_27.INJECT1_1 = "NO";
    CCU2D add_33919_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48158), .COUT(n48159));
    defparam add_33919_25.INIT0 = 16'hf555;
    defparam add_33919_25.INIT1 = 16'hf555;
    defparam add_33919_25.INJECT1_0 = "NO";
    defparam add_33919_25.INJECT1_1 = "NO";
    CCU2D add_33919_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48157), .COUT(n48158));
    defparam add_33919_23.INIT0 = 16'hf555;
    defparam add_33919_23.INIT1 = 16'hf555;
    defparam add_33919_23.INJECT1_0 = "NO";
    defparam add_33919_23.INJECT1_1 = "NO";
    CCU2D add_33919_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48156), .COUT(n48157));
    defparam add_33919_21.INIT0 = 16'hf555;
    defparam add_33919_21.INIT1 = 16'hf555;
    defparam add_33919_21.INJECT1_0 = "NO";
    defparam add_33919_21.INJECT1_1 = "NO";
    CCU2D add_33919_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48155), .COUT(n48156));
    defparam add_33919_19.INIT0 = 16'hf555;
    defparam add_33919_19.INIT1 = 16'hf555;
    defparam add_33919_19.INJECT1_0 = "NO";
    defparam add_33919_19.INJECT1_1 = "NO";
    CCU2D add_33919_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48154), .COUT(n48155));
    defparam add_33919_17.INIT0 = 16'hf555;
    defparam add_33919_17.INIT1 = 16'hf555;
    defparam add_33919_17.INJECT1_0 = "NO";
    defparam add_33919_17.INJECT1_1 = "NO";
    CCU2D add_33919_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48153), .COUT(n48154));
    defparam add_33919_15.INIT0 = 16'hf555;
    defparam add_33919_15.INIT1 = 16'hf555;
    defparam add_33919_15.INJECT1_0 = "NO";
    defparam add_33919_15.INJECT1_1 = "NO";
    CCU2D add_33919_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48152), .COUT(n48153));
    defparam add_33919_13.INIT0 = 16'hf555;
    defparam add_33919_13.INIT1 = 16'hf555;
    defparam add_33919_13.INJECT1_0 = "NO";
    defparam add_33919_13.INJECT1_1 = "NO";
    CCU2D add_33919_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48151), .COUT(n48152));
    defparam add_33919_11.INIT0 = 16'hf555;
    defparam add_33919_11.INIT1 = 16'hf555;
    defparam add_33919_11.INJECT1_0 = "NO";
    defparam add_33919_11.INJECT1_1 = "NO";
    CCU2D add_33919_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48150), .COUT(n48151));
    defparam add_33919_9.INIT0 = 16'hf555;
    defparam add_33919_9.INIT1 = 16'hf555;
    defparam add_33919_9.INJECT1_0 = "NO";
    defparam add_33919_9.INJECT1_1 = "NO";
    CCU2D add_33919_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48149), .COUT(n48150));
    defparam add_33919_7.INIT0 = 16'hf555;
    defparam add_33919_7.INIT1 = 16'hf555;
    defparam add_33919_7.INJECT1_0 = "NO";
    defparam add_33919_7.INJECT1_1 = "NO";
    CCU2D add_33919_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48148), .COUT(n48149));
    defparam add_33919_5.INIT0 = 16'hf555;
    defparam add_33919_5.INIT1 = 16'hf555;
    defparam add_33919_5.INJECT1_0 = "NO";
    defparam add_33919_5.INJECT1_1 = "NO";
    CCU2D add_33919_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48147), .COUT(n48148));
    defparam add_33919_3.INIT0 = 16'hf555;
    defparam add_33919_3.INIT1 = 16'hf555;
    defparam add_33919_3.INJECT1_0 = "NO";
    defparam add_33919_3.INJECT1_1 = "NO";
    CCU2D add_33919_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48147));
    defparam add_33919_1.INIT0 = 16'hF000;
    defparam add_33919_1.INIT1 = 16'ha666;
    defparam add_33919_1.INJECT1_0 = "NO";
    defparam add_33919_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54619), .C(n13241), .D(n54825), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    LUT4 mux_2052_i2_4_lut (.A(n68), .B(n15006[0]), .C(n6831), .D(n52733), 
         .Z(n6832[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2052_i4_4_lut (.A(n39343), .B(n54724), .C(n6831), .D(n4), 
         .Z(n6832[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42588), .B(n54556), .C(n447[3]), .D(n54684), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2052_i8_4_lut (.A(n6656[7]), .B(n54724), .C(n6831), .D(n54556), 
         .Z(n6832[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i8_4_lut.init = 16'h303a;
    LUT4 mux_2052_i9_4_lut (.A(n6656[8]), .B(n54724), .C(n6831), .D(n54556), 
         .Z(n6832[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i9_4_lut.init = 16'h303a;
    LUT4 mux_2052_i10_4_lut (.A(n76), .B(n54724), .C(n6831), .D(n54556), 
         .Z(n6832[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i10_4_lut.init = 16'h303a;
    LUT4 mux_2052_i13_4_lut (.A(n54556), .B(n54724), .C(n6831), .D(n103), 
         .Z(n6832[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2052_i13_4_lut.init = 16'h3530;
    LUT4 i1_2_lut_rep_616 (.A(n42588), .B(n13206), .Z(n54619)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_616.init = 16'h8888;
    LUT4 i1_2_lut_rep_604_3_lut (.A(n42588), .B(n13206), .C(state[1]), 
         .Z(n54607)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_604_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42588), .B(n13206), .C(n54684), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    CCU2D add_3112_33 (.A0(bit_counter[31]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48338), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_33.INIT0 = 16'h5999;
    defparam add_3112_33.INIT1 = 16'h0000;
    defparam add_3112_33.INJECT1_0 = "NO";
    defparam add_3112_33.INJECT1_1 = "NO";
    CCU2D add_3112_31 (.A0(bit_counter[29]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48337), .COUT(n48338), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_31.INIT0 = 16'h5999;
    defparam add_3112_31.INIT1 = 16'h5999;
    defparam add_3112_31.INJECT1_0 = "NO";
    defparam add_3112_31.INJECT1_1 = "NO";
    CCU2D add_3112_29 (.A0(bit_counter[27]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48336), .COUT(n48337), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_29.INIT0 = 16'h5999;
    defparam add_3112_29.INIT1 = 16'h5999;
    defparam add_3112_29.INJECT1_0 = "NO";
    defparam add_3112_29.INJECT1_1 = "NO";
    CCU2D add_3112_27 (.A0(bit_counter[25]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48335), .COUT(n48336), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_27.INIT0 = 16'h5999;
    defparam add_3112_27.INIT1 = 16'h5999;
    defparam add_3112_27.INJECT1_0 = "NO";
    defparam add_3112_27.INJECT1_1 = "NO";
    CCU2D add_3112_25 (.A0(bit_counter[23]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48334), .COUT(n48335), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_25.INIT0 = 16'h5999;
    defparam add_3112_25.INIT1 = 16'h5999;
    defparam add_3112_25.INJECT1_0 = "NO";
    defparam add_3112_25.INJECT1_1 = "NO";
    CCU2D add_3112_23 (.A0(bit_counter[21]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48333), .COUT(n48334), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_23.INIT0 = 16'h5999;
    defparam add_3112_23.INIT1 = 16'h5999;
    defparam add_3112_23.INJECT1_0 = "NO";
    defparam add_3112_23.INJECT1_1 = "NO";
    CCU2D add_3112_21 (.A0(bit_counter[19]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48332), .COUT(n48333), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_21.INIT0 = 16'h5999;
    defparam add_3112_21.INIT1 = 16'h5999;
    defparam add_3112_21.INJECT1_0 = "NO";
    defparam add_3112_21.INJECT1_1 = "NO";
    CCU2D add_3112_19 (.A0(bit_counter[17]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48331), .COUT(n48332), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_19.INIT0 = 16'h5999;
    defparam add_3112_19.INIT1 = 16'h5999;
    defparam add_3112_19.INJECT1_0 = "NO";
    defparam add_3112_19.INJECT1_1 = "NO";
    CCU2D add_3112_17 (.A0(bit_counter[15]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48330), .COUT(n48331), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_17.INIT0 = 16'h5999;
    defparam add_3112_17.INIT1 = 16'h5999;
    defparam add_3112_17.INJECT1_0 = "NO";
    defparam add_3112_17.INJECT1_1 = "NO";
    CCU2D add_3112_15 (.A0(bit_counter[13]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48329), .COUT(n48330), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_15.INIT0 = 16'h5999;
    defparam add_3112_15.INIT1 = 16'h5999;
    defparam add_3112_15.INJECT1_0 = "NO";
    defparam add_3112_15.INJECT1_1 = "NO";
    CCU2D add_3112_13 (.A0(bit_counter[11]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48328), .COUT(n48329), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_13.INIT0 = 16'h5999;
    defparam add_3112_13.INIT1 = 16'h5999;
    defparam add_3112_13.INJECT1_0 = "NO";
    defparam add_3112_13.INJECT1_1 = "NO";
    CCU2D add_3112_11 (.A0(bit_counter[9]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48327), .COUT(n48328), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_11.INIT0 = 16'h5999;
    defparam add_3112_11.INIT1 = 16'h5999;
    defparam add_3112_11.INJECT1_0 = "NO";
    defparam add_3112_11.INJECT1_1 = "NO";
    CCU2D add_3112_9 (.A0(bit_counter[7]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48326), .COUT(n48327), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_9.INIT0 = 16'h5999;
    defparam add_3112_9.INIT1 = 16'h5999;
    defparam add_3112_9.INJECT1_0 = "NO";
    defparam add_3112_9.INJECT1_1 = "NO";
    CCU2D add_3112_7 (.A0(bit_counter[5]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48325), .COUT(n48326), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_7.INIT0 = 16'h5999;
    defparam add_3112_7.INIT1 = 16'h5999;
    defparam add_3112_7.INJECT1_0 = "NO";
    defparam add_3112_7.INJECT1_1 = "NO";
    CCU2D add_3112_5 (.A0(bit_counter[3]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48324), .COUT(n48325), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_5.INIT0 = 16'h5999;
    defparam add_3112_5.INIT1 = 16'h5999;
    defparam add_3112_5.INJECT1_0 = "NO";
    defparam add_3112_5.INJECT1_1 = "NO";
    CCU2D add_3112_3 (.A0(bit_counter[1]), .B0(n13206), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13206), .C1(GND_net), 
          .D1(GND_net), .CIN(n48323), .COUT(n48324), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_3.INIT0 = 16'h5999;
    defparam add_3112_3.INIT1 = 16'h5999;
    defparam add_3112_3.INJECT1_0 = "NO";
    defparam add_3112_3.INJECT1_1 = "NO";
    CCU2D add_3112_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13206), .C1(GND_net), .D1(GND_net), 
          .COUT(n48323), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3112_1.INIT0 = 16'hF000;
    defparam add_3112_1.INIT1 = 16'h5999;
    defparam add_3112_1.INJECT1_0 = "NO";
    defparam add_3112_1.INJECT1_1 = "NO";
    PFUMX i38961 (.BLUT(n54980), .ALUT(n54981), .C0(state[0]), .Z(n54982));
    PFUMX i38923 (.BLUT(n54922), .ALUT(n54923), .C0(state[1]), .Z(n54924));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U24 
//

module \WS2812(48000000,"111111111")_U24  (sclk_c, \port_status[4] , ws2813_out_c_4, 
            \Q[4] , \RdAddress[4] , GND_net);
    input sclk_c;
    output \port_status[4] ;
    output ws2813_out_c_4;
    input [23:0]\Q[4] ;
    output [8:0]\RdAddress[4] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_905;
    wire [31:0]n7144;
    
    wire sclk_c_enable_43, n54818, sclk_c_enable_44, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_47;
    wire [2:0]state_2__N_104;
    wire [31:0]n447;
    
    wire n13171, n54911, n13136, n54910, n54938, n42592, n55531, 
        n54937, n54965, n54964, n54599, n54990, n54989, n54715;
    wire [31:0]n6968;
    
    wire n54654, n23, n54716, n25, n53268, n53269;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53270, n34936, sclk_c_enable_1206, n42538;
    wire [6:0]n15014;
    
    wire sclk_c_enable_1205;
    wire [31:0]bit_counter_31__N_204;
    wire [31:0]bit_counter_31__N_172;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n54798;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1207, n1, n1_adj_908, n34940;
    wire [31:0]n7070;
    
    wire n54912, serial_N_437, n52981, n52982, n52989, n52983, n52984, 
        n52990, n52985, n52986, n52991, n52987, n52988, n52992;
    wire [8:0]n118;
    
    wire n52995, n54884, n53267, n53266, n53265, n53264, n54883, 
        n52993, n52994, n47650, n47649, n47648, n47647, n47646, 
        n47645, n47644, n52673, n15, n14, n47643, n47642, n47641, 
        n47640, n49070, n49069, n49068, n49067, n47639, n49066, 
        n47638, n49065, n49064, n49063, n49062, n49061, n49060, 
        n49059, n49058, n49057, n49056, n49055, n47637, n49007, 
        n49006, n49005, n49004, n49003, n49002, n49001, n49000, 
        n48999, n48998, n48997, n48996, n48995, n48994, n48993, 
        n48992, n47636, n47635, n47617, n47616, n47615, n47614, 
        n48354, n48353, n48352, n48351, n48350, n48349, n48348, 
        n48347, n48346, n48345, n48344, n48343, n48342, n48341, 
        n48340, n48339;
    
    FD1P3AX delay_counter_i0_i0 (.D(n7144[0]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54818), .SP(sclk_c_enable_43), .CK(sclk_c), 
            .Q(\port_status[4] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_44), .CK(sclk_c), 
            .Q(ws2813_out_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_47), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_47), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_47), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 mux_2126_i3_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13171), .Z(n54911)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2126_i3_4_lut_then_4_lut.init = 16'hb1f0;
    LUT4 mux_2126_i3_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13136), .Z(n54910)) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2126_i3_4_lut_else_4_lut.init = 16'hb0f4;
    LUT4 i1_3_lut_4_lut_4_lut_then_2_lut (.A(n13171), .B(state[2]), .Z(n54938)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_3_lut_4_lut_4_lut_then_2_lut.init = 16'h2222;
    LUT4 i29244_2_lut_rep_842 (.A(n42592), .B(n13136), .Z(n55531)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29244_2_lut_rep_842.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut_else_2_lut_4_lut (.A(n42592), .B(n13136), 
         .C(state[0]), .D(state[2]), .Z(n54937)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_else_2_lut_4_lut.init = 16'h0070;
    LUT4 mux_2821_i3_then_3_lut (.A(state[2]), .B(state[0]), .C(n13171), 
         .Z(n54965)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam mux_2821_i3_then_3_lut.init = 16'h4040;
    LUT4 mux_2821_i3_else_3_lut (.A(state[2]), .B(state[0]), .C(n42592), 
         .D(n13136), .Z(n54964)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam mux_2821_i3_else_3_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_596_3_lut (.A(state[2]), .B(n13171), .C(state[1]), 
         .Z(n54599)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_596_3_lut.init = 16'h4040;
    LUT4 mux_2821_i1_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(n13171), .Z(n54990)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B (C (D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2821_i1_4_lut_then_4_lut.init = 16'h175f;
    LUT4 mux_2821_i1_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(n13171), .Z(n54989)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B ((D)+!C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2821_i1_4_lut_else_4_lut.init = 16'h135b;
    LUT4 mux_2120_i8_3_lut_4_lut (.A(n42592), .B(n13136), .C(n54715), 
         .D(n447[7]), .Z(n6968[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2120_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2120_i9_3_lut_4_lut (.A(n42592), .B(n13136), .C(n54715), 
         .D(n447[8]), .Z(n6968[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2120_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2120_i10_3_lut_4_lut (.A(n42592), .B(n13136), .C(n54715), 
         .D(n447[9]), .Z(n6968[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2120_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2120_i13_3_lut_4_lut (.A(n42592), .B(n13136), .C(n54715), 
         .D(n447[12]), .Z(n6968[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2120_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i2148_3_lut_rep_651 (.A(state[2]), .B(state[1]), .C(n13171), 
         .Z(n54654)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2148_3_lut_rep_651.init = 16'ha8a8;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(n447[0]), 
         .D(state[0]), .Z(n23)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i2_2_lut_rep_713_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54716)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2_2_lut_rep_713_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_502 (.A(state[2]), .B(state[1]), .C(n447[1]), 
         .D(state[0]), .Z(n25)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_502.init = 16'he0f0;
    L6MUX21 i38064 (.D0(n53268), .D1(n53269), .SD(bit_counter[2]), .Z(n53270));
    LUT4 i38615_2_lut_rep_549_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(n13171), .D(state[2]), .Z(sclk_c_enable_905)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i38615_2_lut_rep_549_2_lut_3_lut_4_lut.init = 16'hffef;
    LUT4 i22724_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut (.A(state[1]), .B(n13171), 
         .C(state[2]), .Z(n34936)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i22724_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut.init = 16'he0e0;
    LUT4 i27326_3_lut_3_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(sclk_c_enable_1206)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam i27326_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i30369_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42538)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i30369_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i28675_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15014[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28675_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13171), 
         .Z(sclk_c_enable_44)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_rep_712_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .Z(n54715)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_712_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13136), 
         .D(state[1]), .Z(sclk_c_enable_1205)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i37709_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13171), 
         .D(state[1]), .Z(sclk_c_enable_47)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i37709_3_lut_4_lut_4_lut_4_lut.init = 16'hfcf2;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_503 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_503.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_504 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_504.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_505 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_505.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_506 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_506.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_507 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_507.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_508 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_508.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_509 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_509.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_510 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_510.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_511 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_511.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_512 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_512.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_513 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_513.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_514 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_514.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_515 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_515.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_516 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_516.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_517 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_517.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_518 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_518.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_519 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_519.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_520 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_520.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_521 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_521.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_522 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_522.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_523 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_523.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_524 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_524.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_525 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_525.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_526 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_526.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_527 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_527.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_528 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_528.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_529 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_529.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_530 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_530.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_531 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_531.init = 16'h2020;
    FD1P3IX pixel_i23 (.D(\Q[4] [23]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[4] [22]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[4] [21]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[4] [20]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[4] [19]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[4] [18]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[4] [17]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[4] [16]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[4] [15]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[4] [14]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[4] [13]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[4] [12]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[4] [11]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[4] [10]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[4] [9]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[4] [8]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[4] [7]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[4] [6]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[4] [5]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[4] [4]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[4] [3]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[4] [2]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[4] [1]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1207), .CD(n54798), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_908), .SP(sclk_c_enable_1207), .CD(n54798), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_905), 
            .CD(n34940), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_905), .CD(n34940), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_905), .CD(n34940), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n7070[4]), .SP(sclk_c_enable_905), .CD(n34936), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54912), .SP(sclk_c_enable_905), .CD(n34936), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i38416_2_lut_rep_803 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1207)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38416_2_lut_rep_803.init = 16'h9999;
    LUT4 i22877_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n54798)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22877_2_lut_2_lut.init = 16'h8888;
    FD1P3AX delay_counter_i0_i1 (.D(n7144[1]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n7144[3]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n7144[7]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n7144[8]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n7144[9]), .SP(sclk_c_enable_905), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n7144[12]), .SP(sclk_c_enable_905), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i27314_1_lut_rep_815 (.A(state[2]), .Z(n54818)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27314_1_lut_rep_815.init = 16'h5555;
    LUT4 i28869_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28869_3_lut_3_lut.init = 16'h5151;
    PFUMX i37783 (.BLUT(n52981), .ALUT(n52982), .C0(bit_counter[1]), .Z(n52989));
    PFUMX i37784 (.BLUT(n52983), .ALUT(n52984), .C0(bit_counter[1]), .Z(n52990));
    PFUMX i37785 (.BLUT(n52985), .ALUT(n52986), .C0(bit_counter[1]), .Z(n52991));
    PFUMX i37786 (.BLUT(n52987), .ALUT(n52988), .C0(bit_counter[1]), .Z(n52992));
    FD1P3IX pixel_i0 (.D(\Q[4] [0]), .SP(sclk_c_enable_1206), .CD(n54798), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1205), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1206), 
            .CD(n54798), .CK(sclk_c), .Q(\RdAddress[4] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1207), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=179, LSE_RLINE=179 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_532 (.A(state[2]), .B(n42592), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_532.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_533 (.A(state[2]), .B(n42592), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_533.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_534 (.A(state[2]), .B(n42592), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_534.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_535 (.A(state[2]), .B(n42592), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_535.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_536 (.A(state[2]), .B(n42592), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_536.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_537 (.A(state[2]), .B(n42592), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_537.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_538 (.A(state[2]), .B(n42592), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_538.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_539 (.A(state[2]), .B(n42592), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_539.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_540 (.A(state[2]), .B(n42592), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_540.init = 16'h1010;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n52995), .B(n53270), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2821_i2_3_lut_4_lut_then_3_lut (.A(state[1]), .B(state[2]), 
         .C(n13136), .Z(n54884)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam mux_2821_i2_3_lut_4_lut_then_3_lut.init = 16'h0101;
    LUT4 i38061_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38061_3_lut.init = 16'hcaca;
    LUT4 i38060_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38060_3_lut.init = 16'hcaca;
    LUT4 i38059_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38059_3_lut.init = 16'hcaca;
    LUT4 i38058_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38058_3_lut.init = 16'hcaca;
    LUT4 mux_2821_i2_3_lut_4_lut_else_3_lut (.A(state[1]), .B(state[2]), 
         .C(n13171), .Z(n54883)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam mux_2821_i2_3_lut_4_lut_else_3_lut.init = 16'h2020;
    LUT4 i28693_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28693_2_lut.init = 16'hbbbb;
    LUT4 i28694_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_908)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28694_2_lut.init = 16'hbbbb;
    L6MUX21 i37789 (.D0(n52993), .D1(n52994), .SD(bit_counter[3]), .Z(n52995));
    PFUMX i38897 (.BLUT(n54883), .ALUT(n54884), .C0(state[0]), .Z(state_2__N_104[1]));
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47650), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47649), .COUT(n47650), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47648), .COUT(n47649), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47647), .COUT(n47648), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    PFUMX i38062 (.BLUT(n53264), .ALUT(n53265), .C0(bit_counter[1]), .Z(n53268));
    PFUMX i38063 (.BLUT(n53266), .ALUT(n53267), .C0(bit_counter[1]), .Z(n53269));
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47646), .COUT(n47647), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47645), .COUT(n47646), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47644), .COUT(n47645), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    LUT4 mux_2136_i1_4_lut (.A(n23), .B(n15014[0]), .C(n54654), .D(n52673), 
         .Z(n7144[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i1_4_lut.init = 16'hcfca;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[3]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42592)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[4]), .C(cur_pixel[2]), 
         .D(cur_pixel[8]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[7]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47643), .COUT(n47644), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47642), .COUT(n47643), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47641), .COUT(n47642), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    LUT4 i22748_4_lut (.A(sclk_c_enable_905), .B(n54599), .C(n54654), 
         .D(n54715), .Z(n34940)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22748_4_lut.init = 16'haaa8;
    LUT4 mux_2126_i5_4_lut (.A(n447[4]), .B(state[0]), .C(n54599), .D(n54715), 
         .Z(n7070[4])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2126_i5_4_lut.init = 16'hc0ca;
    L6MUX21 i37787 (.D0(n52989), .D1(n52990), .SD(bit_counter[2]), .Z(n52993));
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47640), .COUT(n47641), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    L6MUX21 i37788 (.D0(n52991), .D1(n52992), .SD(bit_counter[2]), .Z(n52994));
    CCU2D add_33924_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49070), 
          .S0(n13171));
    defparam add_33924_cout.INIT0 = 16'h0000;
    defparam add_33924_cout.INIT1 = 16'h0000;
    defparam add_33924_cout.INJECT1_0 = "NO";
    defparam add_33924_cout.INJECT1_1 = "NO";
    CCU2D add_33924_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49069), .COUT(n49070));
    defparam add_33924_31.INIT0 = 16'hf555;
    defparam add_33924_31.INIT1 = 16'h5555;
    defparam add_33924_31.INJECT1_0 = "NO";
    defparam add_33924_31.INJECT1_1 = "NO";
    CCU2D add_33924_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49068), .COUT(n49069));
    defparam add_33924_29.INIT0 = 16'hf555;
    defparam add_33924_29.INIT1 = 16'hf555;
    defparam add_33924_29.INJECT1_0 = "NO";
    defparam add_33924_29.INJECT1_1 = "NO";
    CCU2D add_33924_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49067), .COUT(n49068));
    defparam add_33924_27.INIT0 = 16'hf555;
    defparam add_33924_27.INIT1 = 16'hf555;
    defparam add_33924_27.INJECT1_0 = "NO";
    defparam add_33924_27.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47639), .COUT(n47640), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_33924_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49066), .COUT(n49067));
    defparam add_33924_25.INIT0 = 16'hf555;
    defparam add_33924_25.INIT1 = 16'hf555;
    defparam add_33924_25.INJECT1_0 = "NO";
    defparam add_33924_25.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47638), .COUT(n47639), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_33924_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49065), .COUT(n49066));
    defparam add_33924_23.INIT0 = 16'hf555;
    defparam add_33924_23.INIT1 = 16'hf555;
    defparam add_33924_23.INJECT1_0 = "NO";
    defparam add_33924_23.INJECT1_1 = "NO";
    CCU2D add_33924_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49064), .COUT(n49065));
    defparam add_33924_21.INIT0 = 16'hf555;
    defparam add_33924_21.INIT1 = 16'hf555;
    defparam add_33924_21.INJECT1_0 = "NO";
    defparam add_33924_21.INJECT1_1 = "NO";
    CCU2D add_33924_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49063), .COUT(n49064));
    defparam add_33924_19.INIT0 = 16'hf555;
    defparam add_33924_19.INIT1 = 16'hf555;
    defparam add_33924_19.INJECT1_0 = "NO";
    defparam add_33924_19.INJECT1_1 = "NO";
    CCU2D add_33924_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49062), .COUT(n49063));
    defparam add_33924_17.INIT0 = 16'hf555;
    defparam add_33924_17.INIT1 = 16'hf555;
    defparam add_33924_17.INJECT1_0 = "NO";
    defparam add_33924_17.INJECT1_1 = "NO";
    CCU2D add_33924_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49061), .COUT(n49062));
    defparam add_33924_15.INIT0 = 16'hf555;
    defparam add_33924_15.INIT1 = 16'hf555;
    defparam add_33924_15.INJECT1_0 = "NO";
    defparam add_33924_15.INJECT1_1 = "NO";
    CCU2D add_33924_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49060), .COUT(n49061));
    defparam add_33924_13.INIT0 = 16'hf555;
    defparam add_33924_13.INIT1 = 16'hf555;
    defparam add_33924_13.INJECT1_0 = "NO";
    defparam add_33924_13.INJECT1_1 = "NO";
    CCU2D add_33924_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49059), .COUT(n49060));
    defparam add_33924_11.INIT0 = 16'hf555;
    defparam add_33924_11.INIT1 = 16'hf555;
    defparam add_33924_11.INJECT1_0 = "NO";
    defparam add_33924_11.INJECT1_1 = "NO";
    CCU2D add_33924_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49058), .COUT(n49059));
    defparam add_33924_9.INIT0 = 16'hf555;
    defparam add_33924_9.INIT1 = 16'hf555;
    defparam add_33924_9.INJECT1_0 = "NO";
    defparam add_33924_9.INJECT1_1 = "NO";
    CCU2D add_33924_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49057), .COUT(n49058));
    defparam add_33924_7.INIT0 = 16'hf555;
    defparam add_33924_7.INIT1 = 16'hf555;
    defparam add_33924_7.INJECT1_0 = "NO";
    defparam add_33924_7.INJECT1_1 = "NO";
    CCU2D add_33924_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49056), .COUT(n49057));
    defparam add_33924_5.INIT0 = 16'hf555;
    defparam add_33924_5.INIT1 = 16'hf555;
    defparam add_33924_5.INJECT1_0 = "NO";
    defparam add_33924_5.INJECT1_1 = "NO";
    CCU2D add_33924_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49055), .COUT(n49056));
    defparam add_33924_3.INIT0 = 16'hf555;
    defparam add_33924_3.INIT1 = 16'hf555;
    defparam add_33924_3.INJECT1_0 = "NO";
    defparam add_33924_3.INJECT1_1 = "NO";
    CCU2D add_33924_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n49055));
    defparam add_33924_1.INIT0 = 16'hF000;
    defparam add_33924_1.INIT1 = 16'ha666;
    defparam add_33924_1.INJECT1_0 = "NO";
    defparam add_33924_1.INJECT1_1 = "NO";
    LUT4 i37782_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n52988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37782_3_lut.init = 16'hcaca;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47637), .COUT(n47638), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_33926_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49007), 
          .S0(n13136));
    defparam add_33926_cout.INIT0 = 16'h0000;
    defparam add_33926_cout.INIT1 = 16'h0000;
    defparam add_33926_cout.INJECT1_0 = "NO";
    defparam add_33926_cout.INJECT1_1 = "NO";
    CCU2D add_33926_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49006), .COUT(n49007));
    defparam add_33926_31.INIT0 = 16'hf555;
    defparam add_33926_31.INIT1 = 16'h5555;
    defparam add_33926_31.INJECT1_0 = "NO";
    defparam add_33926_31.INJECT1_1 = "NO";
    LUT4 i37781_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n52987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37781_3_lut.init = 16'hcaca;
    CCU2D add_33926_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49005), .COUT(n49006));
    defparam add_33926_29.INIT0 = 16'hf555;
    defparam add_33926_29.INIT1 = 16'hf555;
    defparam add_33926_29.INJECT1_0 = "NO";
    defparam add_33926_29.INJECT1_1 = "NO";
    CCU2D add_33926_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49004), .COUT(n49005));
    defparam add_33926_27.INIT0 = 16'hf555;
    defparam add_33926_27.INIT1 = 16'hf555;
    defparam add_33926_27.INJECT1_0 = "NO";
    defparam add_33926_27.INJECT1_1 = "NO";
    CCU2D add_33926_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49003), .COUT(n49004));
    defparam add_33926_25.INIT0 = 16'hf555;
    defparam add_33926_25.INIT1 = 16'hf555;
    defparam add_33926_25.INJECT1_0 = "NO";
    defparam add_33926_25.INJECT1_1 = "NO";
    LUT4 i37780_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n52986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37780_3_lut.init = 16'hcaca;
    LUT4 i37779_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n52985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37779_3_lut.init = 16'hcaca;
    CCU2D add_33926_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49002), .COUT(n49003));
    defparam add_33926_23.INIT0 = 16'hf555;
    defparam add_33926_23.INIT1 = 16'hf555;
    defparam add_33926_23.INJECT1_0 = "NO";
    defparam add_33926_23.INJECT1_1 = "NO";
    CCU2D add_33926_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49001), .COUT(n49002));
    defparam add_33926_21.INIT0 = 16'hf555;
    defparam add_33926_21.INIT1 = 16'hf555;
    defparam add_33926_21.INJECT1_0 = "NO";
    defparam add_33926_21.INJECT1_1 = "NO";
    CCU2D add_33926_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49000), .COUT(n49001));
    defparam add_33926_19.INIT0 = 16'hf555;
    defparam add_33926_19.INIT1 = 16'hf555;
    defparam add_33926_19.INJECT1_0 = "NO";
    defparam add_33926_19.INJECT1_1 = "NO";
    CCU2D add_33926_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48999), .COUT(n49000));
    defparam add_33926_17.INIT0 = 16'hf555;
    defparam add_33926_17.INIT1 = 16'hf555;
    defparam add_33926_17.INJECT1_0 = "NO";
    defparam add_33926_17.INJECT1_1 = "NO";
    CCU2D add_33926_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48998), .COUT(n48999));
    defparam add_33926_15.INIT0 = 16'hf555;
    defparam add_33926_15.INIT1 = 16'hf555;
    defparam add_33926_15.INJECT1_0 = "NO";
    defparam add_33926_15.INJECT1_1 = "NO";
    CCU2D add_33926_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48997), .COUT(n48998));
    defparam add_33926_13.INIT0 = 16'hf555;
    defparam add_33926_13.INIT1 = 16'hf555;
    defparam add_33926_13.INJECT1_0 = "NO";
    defparam add_33926_13.INJECT1_1 = "NO";
    CCU2D add_33926_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48996), .COUT(n48997));
    defparam add_33926_11.INIT0 = 16'hf555;
    defparam add_33926_11.INIT1 = 16'hf555;
    defparam add_33926_11.INJECT1_0 = "NO";
    defparam add_33926_11.INJECT1_1 = "NO";
    CCU2D add_33926_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48995), .COUT(n48996));
    defparam add_33926_9.INIT0 = 16'hf555;
    defparam add_33926_9.INIT1 = 16'hf555;
    defparam add_33926_9.INJECT1_0 = "NO";
    defparam add_33926_9.INJECT1_1 = "NO";
    CCU2D add_33926_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48994), .COUT(n48995));
    defparam add_33926_7.INIT0 = 16'hf555;
    defparam add_33926_7.INIT1 = 16'hf555;
    defparam add_33926_7.INJECT1_0 = "NO";
    defparam add_33926_7.INJECT1_1 = "NO";
    CCU2D add_33926_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48993), .COUT(n48994));
    defparam add_33926_5.INIT0 = 16'hf555;
    defparam add_33926_5.INIT1 = 16'hf555;
    defparam add_33926_5.INJECT1_0 = "NO";
    defparam add_33926_5.INJECT1_1 = "NO";
    CCU2D add_33926_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48992), .COUT(n48993));
    defparam add_33926_3.INIT0 = 16'hf555;
    defparam add_33926_3.INIT1 = 16'hf555;
    defparam add_33926_3.INJECT1_0 = "NO";
    defparam add_33926_3.INJECT1_1 = "NO";
    CCU2D add_33926_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48992));
    defparam add_33926_1.INIT0 = 16'hF000;
    defparam add_33926_1.INIT1 = 16'ha666;
    defparam add_33926_1.INJECT1_0 = "NO";
    defparam add_33926_1.INJECT1_1 = "NO";
    LUT4 i37778_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37778_3_lut.init = 16'hcaca;
    LUT4 i37777_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37777_3_lut.init = 16'hcaca;
    LUT4 i37776_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37776_3_lut.init = 16'hcaca;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47636), .COUT(n47637), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47635), .COUT(n47636), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47635), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i37775_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37775_3_lut.init = 16'hcaca;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47617), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47616), .COUT(n47617), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47615), .COUT(n47616), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    LUT4 mux_2136_i2_4_lut (.A(n25), .B(n15014[0]), .C(n54654), .D(n52673), 
         .Z(n7144[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2136_i4_4_lut (.A(n6968[3]), .B(n42538), .C(n54654), .D(n54599), 
         .Z(n7144[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i4_4_lut.init = 16'h3f3a;
    LUT4 i29592_4_lut (.A(n42592), .B(n447[3]), .C(n54716), .D(n13136), 
         .Z(n6968[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29592_4_lut.init = 16'hcacf;
    LUT4 mux_2136_i8_4_lut (.A(n6968[7]), .B(n42538), .C(n54654), .D(n54599), 
         .Z(n7144[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i8_4_lut.init = 16'h303a;
    LUT4 mux_2136_i9_4_lut (.A(n6968[8]), .B(n42538), .C(n54654), .D(n54599), 
         .Z(n7144[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i9_4_lut.init = 16'h303a;
    LUT4 mux_2136_i10_4_lut (.A(n6968[9]), .B(n42538), .C(n54654), .D(n54599), 
         .Z(n7144[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i10_4_lut.init = 16'h303a;
    LUT4 mux_2136_i13_4_lut (.A(n6968[12]), .B(n42538), .C(n54654), .D(n54599), 
         .Z(n7144[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2136_i13_4_lut.init = 16'h303a;
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47614), .COUT(n47615), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47614), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3110_33 (.A0(bit_counter[31]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48354), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_33.INIT0 = 16'h5999;
    defparam add_3110_33.INIT1 = 16'h0000;
    defparam add_3110_33.INJECT1_0 = "NO";
    defparam add_3110_33.INJECT1_1 = "NO";
    CCU2D add_3110_31 (.A0(bit_counter[29]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48353), .COUT(n48354), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_31.INIT0 = 16'h5999;
    defparam add_3110_31.INIT1 = 16'h5999;
    defparam add_3110_31.INJECT1_0 = "NO";
    defparam add_3110_31.INJECT1_1 = "NO";
    CCU2D add_3110_29 (.A0(bit_counter[27]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48352), .COUT(n48353), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_29.INIT0 = 16'h5999;
    defparam add_3110_29.INIT1 = 16'h5999;
    defparam add_3110_29.INJECT1_0 = "NO";
    defparam add_3110_29.INJECT1_1 = "NO";
    CCU2D add_3110_27 (.A0(bit_counter[25]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48351), .COUT(n48352), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_27.INIT0 = 16'h5999;
    defparam add_3110_27.INIT1 = 16'h5999;
    defparam add_3110_27.INJECT1_0 = "NO";
    defparam add_3110_27.INJECT1_1 = "NO";
    CCU2D add_3110_25 (.A0(bit_counter[23]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48350), .COUT(n48351), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_25.INIT0 = 16'h5999;
    defparam add_3110_25.INIT1 = 16'h5999;
    defparam add_3110_25.INJECT1_0 = "NO";
    defparam add_3110_25.INJECT1_1 = "NO";
    CCU2D add_3110_23 (.A0(bit_counter[21]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48349), .COUT(n48350), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_23.INIT0 = 16'h5999;
    defparam add_3110_23.INIT1 = 16'h5999;
    defparam add_3110_23.INJECT1_0 = "NO";
    defparam add_3110_23.INJECT1_1 = "NO";
    CCU2D add_3110_21 (.A0(bit_counter[19]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48348), .COUT(n48349), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_21.INIT0 = 16'h5999;
    defparam add_3110_21.INIT1 = 16'h5999;
    defparam add_3110_21.INJECT1_0 = "NO";
    defparam add_3110_21.INJECT1_1 = "NO";
    CCU2D add_3110_19 (.A0(bit_counter[17]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48347), .COUT(n48348), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_19.INIT0 = 16'h5999;
    defparam add_3110_19.INIT1 = 16'h5999;
    defparam add_3110_19.INJECT1_0 = "NO";
    defparam add_3110_19.INJECT1_1 = "NO";
    CCU2D add_3110_17 (.A0(bit_counter[15]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48346), .COUT(n48347), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_17.INIT0 = 16'h5999;
    defparam add_3110_17.INIT1 = 16'h5999;
    defparam add_3110_17.INJECT1_0 = "NO";
    defparam add_3110_17.INJECT1_1 = "NO";
    CCU2D add_3110_15 (.A0(bit_counter[13]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48345), .COUT(n48346), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_15.INIT0 = 16'h5999;
    defparam add_3110_15.INIT1 = 16'h5999;
    defparam add_3110_15.INJECT1_0 = "NO";
    defparam add_3110_15.INJECT1_1 = "NO";
    CCU2D add_3110_13 (.A0(bit_counter[11]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48344), .COUT(n48345), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_13.INIT0 = 16'h5999;
    defparam add_3110_13.INIT1 = 16'h5999;
    defparam add_3110_13.INJECT1_0 = "NO";
    defparam add_3110_13.INJECT1_1 = "NO";
    CCU2D add_3110_11 (.A0(bit_counter[9]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48343), .COUT(n48344), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_11.INIT0 = 16'h5999;
    defparam add_3110_11.INIT1 = 16'h5999;
    defparam add_3110_11.INJECT1_0 = "NO";
    defparam add_3110_11.INJECT1_1 = "NO";
    CCU2D add_3110_9 (.A0(bit_counter[7]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48342), .COUT(n48343), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_9.INIT0 = 16'h5999;
    defparam add_3110_9.INIT1 = 16'h5999;
    defparam add_3110_9.INJECT1_0 = "NO";
    defparam add_3110_9.INJECT1_1 = "NO";
    CCU2D add_3110_7 (.A0(bit_counter[5]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48341), .COUT(n48342), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_7.INIT0 = 16'h5999;
    defparam add_3110_7.INIT1 = 16'h5999;
    defparam add_3110_7.INJECT1_0 = "NO";
    defparam add_3110_7.INJECT1_1 = "NO";
    CCU2D add_3110_5 (.A0(bit_counter[3]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48340), .COUT(n48341), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_5.INIT0 = 16'h5999;
    defparam add_3110_5.INIT1 = 16'h5999;
    defparam add_3110_5.INJECT1_0 = "NO";
    defparam add_3110_5.INJECT1_1 = "NO";
    CCU2D add_3110_3 (.A0(bit_counter[1]), .B0(n13136), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13136), .C1(GND_net), 
          .D1(GND_net), .CIN(n48339), .COUT(n48340), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_3.INIT0 = 16'h5999;
    defparam add_3110_3.INIT1 = 16'h5999;
    defparam add_3110_3.INJECT1_0 = "NO";
    defparam add_3110_3.INJECT1_1 = "NO";
    CCU2D add_3110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13136), .C1(GND_net), .D1(GND_net), 
          .COUT(n48339), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3110_1.INIT0 = 16'hF000;
    defparam add_3110_1.INIT1 = 16'h5999;
    defparam add_3110_1.INJECT1_0 = "NO";
    defparam add_3110_1.INJECT1_1 = "NO";
    PFUMX i38967 (.BLUT(n54989), .ALUT(n54990), .C0(n55531), .Z(state_2__N_104[0]));
    PFUMX i38951 (.BLUT(n54964), .ALUT(n54965), .C0(state[1]), .Z(state_2__N_104[2]));
    PFUMX i38933 (.BLUT(n54937), .ALUT(n54938), .C0(state[1]), .Z(n52673));
    PFUMX i38915 (.BLUT(n54910), .ALUT(n54911), .C0(state[1]), .Z(n54912));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U20 
//

module \WS2812(48000000,"111111111")_U20  (GND_net, sclk_c, \port_status[8] , 
            ws2813_out_c_8, \Q[8] , \RdAddress[8] );
    input GND_net;
    input sclk_c;
    output \port_status[8] ;
    output ws2813_out_c_8;
    input [23:0]\Q[8] ;
    output [8:0]\RdAddress[8] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n48295;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n13416;
    wire [31:0]bit_counter_31__N_204;
    
    wire n48296, n48294;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_980;
    wire [31:0]n5854;
    
    wire sclk_c_enable_78, n54807, sclk_c_enable_79, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_82;
    wire [2:0]state_2__N_104;
    
    wire n53049, n53050, n53053, n48293, n48292, n53051, n53052, 
        n53054, n48291, n35320;
    wire [31:0]n447;
    
    wire n35316;
    wire [31:0]n5780;
    
    wire n54997, n13451, n54932, n54931, n54996, n54995, n54658, 
        n54814, n54661, n54660, n54605, n42804, n54602, n53296, 
        n53297, n53298, n54723;
    wire [31:0]n5678;
    
    wire serial_N_437, n80;
    wire [6:0]n14959;
    
    wire n42484, n54813, n71, n35498, sclk_c_enable_2418, n74, n38941, 
        sclk_c_enable_2385;
    wire [31:0]bit_counter_31__N_172;
    
    wire n5853, sclk_c_enable_2449, n35469;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]cur_pixel_8__N_107;
    
    wire n53041, n53042, n53043, n53044, n53045, n53046, n53047, 
        n53048;
    wire [8:0]n118;
    
    wire n52670, n15, n14, n53295, n53294, n53293, n53292, n1, 
        n1_adj_907, n53055;
    wire [2:0]n9340;
    
    wire n9347, n49134, n49133, n49132, n49131, n49130, n49129, 
        n49128, n49127, n49126, n49125, n49124, n49123, n49122, 
        n49121, n49120, n49119, n49118, n49117, n49116, n49115, 
        n49114, n49113, n49112, n49111, n49110, n49109, n49108, 
        n49107, n49106, n49105, n49104, n49103, n47750, n47749, 
        n47748, n47747, n47746, n47745, n47744, n47743, n47742, 
        n47741, n47740, n47739, n47738, n47737, n47736, n47735, 
        n47733, n47732, n47731, n47730, n4, n48306, n48305, n48304, 
        n48303, n48302, n48301, n48300, n48299, n48298, n48297;
    
    CCU2D add_3118_11 (.A0(bit_counter[9]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48295), .COUT(n48296), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_11.INIT0 = 16'h5999;
    defparam add_3118_11.INIT1 = 16'h5999;
    defparam add_3118_11.INJECT1_0 = "NO";
    defparam add_3118_11.INJECT1_1 = "NO";
    CCU2D add_3118_9 (.A0(bit_counter[7]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48294), .COUT(n48295), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_9.INIT0 = 16'h5999;
    defparam add_3118_9.INIT1 = 16'h5999;
    defparam add_3118_9.INJECT1_0 = "NO";
    defparam add_3118_9.INJECT1_1 = "NO";
    FD1P3AX delay_counter_i0_i0 (.D(n5854[0]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54807), .SP(sclk_c_enable_78), .CK(sclk_c), 
            .Q(\port_status[8] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_79), .CK(sclk_c), 
            .Q(ws2813_out_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_82), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_82), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_82), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    L6MUX21 i37847 (.D0(n53049), .D1(n53050), .SD(bit_counter[2]), .Z(n53053));
    CCU2D add_3118_7 (.A0(bit_counter[5]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48293), .COUT(n48294), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_7.INIT0 = 16'h5999;
    defparam add_3118_7.INIT1 = 16'h5999;
    defparam add_3118_7.INJECT1_0 = "NO";
    defparam add_3118_7.INJECT1_1 = "NO";
    CCU2D add_3118_5 (.A0(bit_counter[3]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48292), .COUT(n48293), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_5.INIT0 = 16'h5999;
    defparam add_3118_5.INIT1 = 16'h5999;
    defparam add_3118_5.INJECT1_0 = "NO";
    defparam add_3118_5.INJECT1_1 = "NO";
    L6MUX21 i37848 (.D0(n53051), .D1(n53052), .SD(bit_counter[2]), .Z(n53054));
    CCU2D add_3118_3 (.A0(bit_counter[1]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48291), .COUT(n48292), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_3.INIT0 = 16'h5999;
    defparam add_3118_3.INIT1 = 16'h5999;
    defparam add_3118_3.INJECT1_0 = "NO";
    defparam add_3118_3.INJECT1_1 = "NO";
    CCU2D add_3118_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13416), .C1(GND_net), .D1(GND_net), 
          .COUT(n48291), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_1.INIT0 = 16'hF000;
    defparam add_3118_1.INIT1 = 16'h5999;
    defparam add_3118_1.INJECT1_0 = "NO";
    defparam add_3118_1.INJECT1_1 = "NO";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_980), 
            .CD(n35320), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_980), .CD(n35320), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_980), .CD(n35320), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n5780[4]), .SP(sclk_c_enable_980), .CD(n35316), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54997), .SP(sclk_c_enable_980), .CD(n35316), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13451), .Z(sclk_c_enable_82)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i38627_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n13451), 
         .Z(n54932)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38627_4_lut_then_3_lut.init = 16'h1010;
    LUT4 i38627_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n13416), 
         .Z(n54931)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38627_4_lut_else_3_lut.init = 16'h0404;
    LUT4 mux_1868_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13451), .Z(n54996)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1868_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_1868_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13416), .Z(n54995)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1868_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i1_2_lut_rep_655 (.A(state[1]), .B(n13451), .Z(n54658)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_655.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[1]), .B(n13451), .C(n54814), .D(n54661), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd080;
    LUT4 i1_2_lut_rep_657 (.A(state[2]), .B(n13451), .Z(n54660)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_657.init = 16'h4444;
    LUT4 i1_2_lut_rep_602_3_lut (.A(state[2]), .B(n13451), .C(state[1]), 
         .Z(n54605)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_602_3_lut.init = 16'h4040;
    LUT4 i38598_3_lut_rep_603_4_lut (.A(state[2]), .B(n13451), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_980)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38598_3_lut_rep_603_4_lut.init = 16'hfffb;
    LUT4 i37691_2_lut_rep_658 (.A(n42804), .B(n13416), .Z(n54661)) /* synthesis lut_function=(A (B)) */ ;
    defparam i37691_2_lut_rep_658.init = 16'h8888;
    LUT4 i1_2_lut_rep_599_3_lut (.A(n42804), .B(n13416), .C(state[1]), 
         .Z(n54602)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_599_3_lut.init = 16'h0808;
    L6MUX21 i38092 (.D0(n53296), .D1(n53297), .SD(bit_counter[2]), .Z(n53298));
    LUT4 i1_3_lut_4_lut (.A(n54602), .B(n54814), .C(n447[8]), .D(n54723), 
         .Z(n5678[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i26743_1_lut_rep_804 (.A(state[2]), .Z(n54807)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i26743_1_lut_rep_804.init = 16'h5555;
    LUT4 i28924_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28924_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_3_lut_4_lut_adj_455 (.A(n54602), .B(n54814), .C(n447[12]), 
         .D(n54723), .Z(n5678[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_455.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_456 (.A(n54602), .B(n54814), .C(n447[9]), 
         .D(n54723), .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_456.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_457 (.A(n54602), .B(n54814), .C(n447[7]), 
         .D(n54723), .Z(n5678[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_457.init = 16'hf888;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n14959[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i30315_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42484)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i30315_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_810 (.A(state[1]), .B(state[2]), .Z(n54813)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_810.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_rep_720_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54723)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_720_3_lut.init = 16'hefef;
    LUT4 i23349_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n35498)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i23349_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_725_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_2418)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_725_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut_adj_458 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_458.init = 16'he0f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n13451), 
         .Z(sclk_c_enable_79)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_2_lut_rep_811 (.A(state[2]), .B(state[0]), .Z(n54814)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_811.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_459 (.A(state[2]), .B(state[0]), .C(n13416), 
         .D(state[1]), .Z(n38941)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_459.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13416), 
         .D(state[1]), .Z(sclk_c_enable_2385)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_3_lut_adj_460 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_460.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_461 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_461.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_462 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_462.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_463 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_463.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_464 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_464.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_465 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_465.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_466 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_466.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_467 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_467.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_468 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_468.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_469 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_469.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_470 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_470.init = 16'h4040;
    LUT4 i23128_4_lut (.A(sclk_c_enable_980), .B(n54723), .C(n5853), .D(n54605), 
         .Z(n35320)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23128_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_adj_471 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_471.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_472 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_472.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_473 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_473.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_474 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_474.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_475 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_475.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_476 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_476.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_477 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_477.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_478 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_478.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_479 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_479.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_480 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_480.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_481 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_481.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_482 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_482.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_483 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_483.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_484 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_484.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_485 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_485.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_486 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_486.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_487 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_487.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_488 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_488.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_489 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_489.init = 16'h4040;
    FD1P3AX delay_counter_i0_i1 (.D(n5854[1]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n5854[3]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n5854[7]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n5854[8]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n5854[9]), .SP(sclk_c_enable_980), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n5854[12]), .SP(sclk_c_enable_980), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i38406_2_lut_rep_823 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_2449)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38406_2_lut_rep_823.init = 16'h9999;
    LUT4 i23257_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35469)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23257_2_lut_2_lut.init = 16'h8888;
    FD1P3IX pixel_i0 (.D(\Q[8] [0]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    PFUMX i37843 (.BLUT(n53041), .ALUT(n53042), .C0(bit_counter[1]), .Z(n53049));
    PFUMX i37844 (.BLUT(n53043), .ALUT(n53044), .C0(bit_counter[1]), .Z(n53050));
    PFUMX i37845 (.BLUT(n53045), .ALUT(n53046), .C0(bit_counter[1]), .Z(n53051));
    PFUMX i37846 (.BLUT(n53047), .ALUT(n53048), .C0(bit_counter[1]), .Z(n53052));
    LUT4 i1_2_lut_3_lut_adj_490 (.A(state[2]), .B(n42804), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_490.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_491 (.A(state[2]), .B(n42804), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_491.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_492 (.A(state[2]), .B(n42804), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_492.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_493 (.A(state[2]), .B(n42804), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_493.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_494 (.A(state[2]), .B(n42804), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_494.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_495 (.A(state[2]), .B(n42804), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_495.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_496 (.A(state[2]), .B(n42804), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_496.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_497 (.A(state[2]), .B(n42804), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_497.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_498 (.A(state[2]), .B(n42804), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_498.init = 16'h1010;
    LUT4 mux_1878_i1_4_lut (.A(n74), .B(n14959[0]), .C(n5853), .D(n52670), 
         .Z(n5854[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i1_4_lut.init = 16'hcfca;
    LUT4 i1890_3_lut (.A(state[2]), .B(state[1]), .C(n13451), .Z(n5853)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1890_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[2]), .C(n14), .D(cur_pixel[3]), 
         .Z(n42804)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[1]), .C(cur_pixel[8]), 
         .D(cur_pixel[6]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[4]), .B(cur_pixel[0]), .C(cur_pixel[7]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i38089_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38089_3_lut.init = 16'hcaca;
    LUT4 i38088_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38088_3_lut.init = 16'hcaca;
    LUT4 i38087_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38087_3_lut.init = 16'hcaca;
    LUT4 i38086_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38086_3_lut.init = 16'hcaca;
    LUT4 i28772_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28772_2_lut.init = 16'hbbbb;
    LUT4 i28771_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_907)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28771_2_lut.init = 16'hbbbb;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53055), .B(n53298), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i29515_4_lut (.A(n9340[0]), .B(n9347), .C(state[0]), .D(n54658), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29515_4_lut.init = 16'h0322;
    LUT4 i1_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(n13451), 
         .Z(n9347)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_499 (.A(state[0]), .B(n54813), .C(n13416), 
         .D(n42804), .Z(n9340[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_499.init = 16'hfddd;
    LUT4 mux_1868_i5_4_lut_4_lut (.A(state[0]), .B(n54813), .C(n447[4]), 
         .D(n54605), .Z(n5780[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_1868_i5_4_lut_4_lut.init = 16'haad0;
    LUT4 i1_3_lut_4_lut_4_lut_adj_500 (.A(n54814), .B(state[1]), .C(n54661), 
         .D(n54660), .Z(n52670)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_500.init = 16'hce02;
    L6MUX21 i37849 (.D0(n53053), .D1(n53054), .SD(bit_counter[3]), .Z(n53055));
    LUT4 i37842_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37842_3_lut.init = 16'hcaca;
    LUT4 i37841_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37841_3_lut.init = 16'hcaca;
    LUT4 i37840_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37840_3_lut.init = 16'hcaca;
    LUT4 i37839_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37839_3_lut.init = 16'hcaca;
    LUT4 i37838_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37838_3_lut.init = 16'hcaca;
    LUT4 i37837_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37837_3_lut.init = 16'hcaca;
    PFUMX i38090 (.BLUT(n53292), .ALUT(n53293), .C0(bit_counter[1]), .Z(n53296));
    PFUMX i38091 (.BLUT(n53294), .ALUT(n53295), .C0(bit_counter[1]), .Z(n53297));
    LUT4 i37836_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37836_3_lut.init = 16'hcaca;
    LUT4 i37835_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37835_3_lut.init = 16'hcaca;
    CCU2D add_33920_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49134), 
          .S0(n13451));
    defparam add_33920_cout.INIT0 = 16'h0000;
    defparam add_33920_cout.INIT1 = 16'h0000;
    defparam add_33920_cout.INJECT1_0 = "NO";
    defparam add_33920_cout.INJECT1_1 = "NO";
    CCU2D add_33920_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49133), .COUT(n49134));
    defparam add_33920_31.INIT0 = 16'hf555;
    defparam add_33920_31.INIT1 = 16'h5555;
    defparam add_33920_31.INJECT1_0 = "NO";
    defparam add_33920_31.INJECT1_1 = "NO";
    CCU2D add_33920_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49132), .COUT(n49133));
    defparam add_33920_29.INIT0 = 16'hf555;
    defparam add_33920_29.INIT1 = 16'hf555;
    defparam add_33920_29.INJECT1_0 = "NO";
    defparam add_33920_29.INJECT1_1 = "NO";
    CCU2D add_33920_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49131), .COUT(n49132));
    defparam add_33920_27.INIT0 = 16'hf555;
    defparam add_33920_27.INIT1 = 16'hf555;
    defparam add_33920_27.INJECT1_0 = "NO";
    defparam add_33920_27.INJECT1_1 = "NO";
    CCU2D add_33920_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49130), .COUT(n49131));
    defparam add_33920_25.INIT0 = 16'hf555;
    defparam add_33920_25.INIT1 = 16'hf555;
    defparam add_33920_25.INJECT1_0 = "NO";
    defparam add_33920_25.INJECT1_1 = "NO";
    CCU2D add_33920_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49129), .COUT(n49130));
    defparam add_33920_23.INIT0 = 16'hf555;
    defparam add_33920_23.INIT1 = 16'hf555;
    defparam add_33920_23.INJECT1_0 = "NO";
    defparam add_33920_23.INJECT1_1 = "NO";
    CCU2D add_33920_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49128), .COUT(n49129));
    defparam add_33920_21.INIT0 = 16'hf555;
    defparam add_33920_21.INIT1 = 16'hf555;
    defparam add_33920_21.INJECT1_0 = "NO";
    defparam add_33920_21.INJECT1_1 = "NO";
    CCU2D add_33920_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49127), .COUT(n49128));
    defparam add_33920_19.INIT0 = 16'hf555;
    defparam add_33920_19.INIT1 = 16'hf555;
    defparam add_33920_19.INJECT1_0 = "NO";
    defparam add_33920_19.INJECT1_1 = "NO";
    CCU2D add_33920_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49126), .COUT(n49127));
    defparam add_33920_17.INIT0 = 16'hf555;
    defparam add_33920_17.INIT1 = 16'hf555;
    defparam add_33920_17.INJECT1_0 = "NO";
    defparam add_33920_17.INJECT1_1 = "NO";
    CCU2D add_33920_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49125), .COUT(n49126));
    defparam add_33920_15.INIT0 = 16'hf555;
    defparam add_33920_15.INIT1 = 16'hf555;
    defparam add_33920_15.INJECT1_0 = "NO";
    defparam add_33920_15.INJECT1_1 = "NO";
    CCU2D add_33920_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49124), .COUT(n49125));
    defparam add_33920_13.INIT0 = 16'hf555;
    defparam add_33920_13.INIT1 = 16'hf555;
    defparam add_33920_13.INJECT1_0 = "NO";
    defparam add_33920_13.INJECT1_1 = "NO";
    CCU2D add_33920_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49123), .COUT(n49124));
    defparam add_33920_11.INIT0 = 16'hf555;
    defparam add_33920_11.INIT1 = 16'hf555;
    defparam add_33920_11.INJECT1_0 = "NO";
    defparam add_33920_11.INJECT1_1 = "NO";
    CCU2D add_33920_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49122), .COUT(n49123));
    defparam add_33920_9.INIT0 = 16'hf555;
    defparam add_33920_9.INIT1 = 16'hf555;
    defparam add_33920_9.INJECT1_0 = "NO";
    defparam add_33920_9.INJECT1_1 = "NO";
    CCU2D add_33920_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49121), .COUT(n49122));
    defparam add_33920_7.INIT0 = 16'hf555;
    defparam add_33920_7.INIT1 = 16'hf555;
    defparam add_33920_7.INJECT1_0 = "NO";
    defparam add_33920_7.INJECT1_1 = "NO";
    CCU2D add_33920_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49120), .COUT(n49121));
    defparam add_33920_5.INIT0 = 16'hf555;
    defparam add_33920_5.INIT1 = 16'hf555;
    defparam add_33920_5.INJECT1_0 = "NO";
    defparam add_33920_5.INJECT1_1 = "NO";
    CCU2D add_33920_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49119), .COUT(n49120));
    defparam add_33920_3.INIT0 = 16'hf555;
    defparam add_33920_3.INIT1 = 16'hf555;
    defparam add_33920_3.INJECT1_0 = "NO";
    defparam add_33920_3.INJECT1_1 = "NO";
    CCU2D add_33920_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n49119));
    defparam add_33920_1.INIT0 = 16'hF000;
    defparam add_33920_1.INIT1 = 16'ha666;
    defparam add_33920_1.INJECT1_0 = "NO";
    defparam add_33920_1.INJECT1_1 = "NO";
    CCU2D add_33921_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49118), 
          .S0(n13416));
    defparam add_33921_cout.INIT0 = 16'h0000;
    defparam add_33921_cout.INIT1 = 16'h0000;
    defparam add_33921_cout.INJECT1_0 = "NO";
    defparam add_33921_cout.INJECT1_1 = "NO";
    CCU2D add_33921_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49117), .COUT(n49118));
    defparam add_33921_31.INIT0 = 16'hf555;
    defparam add_33921_31.INIT1 = 16'h5555;
    defparam add_33921_31.INJECT1_0 = "NO";
    defparam add_33921_31.INJECT1_1 = "NO";
    CCU2D add_33921_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49116), .COUT(n49117));
    defparam add_33921_29.INIT0 = 16'hf555;
    defparam add_33921_29.INIT1 = 16'hf555;
    defparam add_33921_29.INJECT1_0 = "NO";
    defparam add_33921_29.INJECT1_1 = "NO";
    CCU2D add_33921_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49115), .COUT(n49116));
    defparam add_33921_27.INIT0 = 16'hf555;
    defparam add_33921_27.INIT1 = 16'hf555;
    defparam add_33921_27.INJECT1_0 = "NO";
    defparam add_33921_27.INJECT1_1 = "NO";
    CCU2D add_33921_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49114), .COUT(n49115));
    defparam add_33921_25.INIT0 = 16'hf555;
    defparam add_33921_25.INIT1 = 16'hf555;
    defparam add_33921_25.INJECT1_0 = "NO";
    defparam add_33921_25.INJECT1_1 = "NO";
    CCU2D add_33921_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49113), .COUT(n49114));
    defparam add_33921_23.INIT0 = 16'hf555;
    defparam add_33921_23.INIT1 = 16'hf555;
    defparam add_33921_23.INJECT1_0 = "NO";
    defparam add_33921_23.INJECT1_1 = "NO";
    CCU2D add_33921_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49112), .COUT(n49113));
    defparam add_33921_21.INIT0 = 16'hf555;
    defparam add_33921_21.INIT1 = 16'hf555;
    defparam add_33921_21.INJECT1_0 = "NO";
    defparam add_33921_21.INJECT1_1 = "NO";
    CCU2D add_33921_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49111), .COUT(n49112));
    defparam add_33921_19.INIT0 = 16'hf555;
    defparam add_33921_19.INIT1 = 16'hf555;
    defparam add_33921_19.INJECT1_0 = "NO";
    defparam add_33921_19.INJECT1_1 = "NO";
    CCU2D add_33921_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49110), .COUT(n49111));
    defparam add_33921_17.INIT0 = 16'hf555;
    defparam add_33921_17.INIT1 = 16'hf555;
    defparam add_33921_17.INJECT1_0 = "NO";
    defparam add_33921_17.INJECT1_1 = "NO";
    CCU2D add_33921_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49109), .COUT(n49110));
    defparam add_33921_15.INIT0 = 16'hf555;
    defparam add_33921_15.INIT1 = 16'hf555;
    defparam add_33921_15.INJECT1_0 = "NO";
    defparam add_33921_15.INJECT1_1 = "NO";
    CCU2D add_33921_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49108), .COUT(n49109));
    defparam add_33921_13.INIT0 = 16'hf555;
    defparam add_33921_13.INIT1 = 16'hf555;
    defparam add_33921_13.INJECT1_0 = "NO";
    defparam add_33921_13.INJECT1_1 = "NO";
    CCU2D add_33921_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49107), .COUT(n49108));
    defparam add_33921_11.INIT0 = 16'hf555;
    defparam add_33921_11.INIT1 = 16'hf555;
    defparam add_33921_11.INJECT1_0 = "NO";
    defparam add_33921_11.INJECT1_1 = "NO";
    CCU2D add_33921_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49106), .COUT(n49107));
    defparam add_33921_9.INIT0 = 16'hf555;
    defparam add_33921_9.INIT1 = 16'hf555;
    defparam add_33921_9.INJECT1_0 = "NO";
    defparam add_33921_9.INJECT1_1 = "NO";
    CCU2D add_33921_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49105), .COUT(n49106));
    defparam add_33921_7.INIT0 = 16'hf555;
    defparam add_33921_7.INIT1 = 16'hf555;
    defparam add_33921_7.INJECT1_0 = "NO";
    defparam add_33921_7.INJECT1_1 = "NO";
    CCU2D add_33921_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49104), .COUT(n49105));
    defparam add_33921_5.INIT0 = 16'hf555;
    defparam add_33921_5.INIT1 = 16'hf555;
    defparam add_33921_5.INJECT1_0 = "NO";
    defparam add_33921_5.INJECT1_1 = "NO";
    CCU2D add_33921_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49103), .COUT(n49104));
    defparam add_33921_3.INIT0 = 16'hf555;
    defparam add_33921_3.INIT1 = 16'hf555;
    defparam add_33921_3.INJECT1_0 = "NO";
    defparam add_33921_3.INJECT1_1 = "NO";
    CCU2D add_33921_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n49103));
    defparam add_33921_1.INIT0 = 16'hF000;
    defparam add_33921_1.INIT1 = 16'ha666;
    defparam add_33921_1.INJECT1_0 = "NO";
    defparam add_33921_1.INJECT1_1 = "NO";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47750), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47749), .COUT(n47750), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47748), .COUT(n47749), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47747), .COUT(n47748), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47746), .COUT(n47747), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47745), .COUT(n47746), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47744), .COUT(n47745), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47743), .COUT(n47744), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47742), .COUT(n47743), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47741), .COUT(n47742), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47740), .COUT(n47741), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47739), .COUT(n47740), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47738), .COUT(n47739), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47737), .COUT(n47738), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47736), .COUT(n47737), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47735), .COUT(n47736), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47735), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47733), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47732), .COUT(n47733), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47731), .COUT(n47732), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47730), .COUT(n47731), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47730), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i23104_2_lut_4_lut (.A(n54660), .B(state[0]), .C(state[1]), .D(n5853), 
         .Z(n35316)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23104_2_lut_4_lut.init = 16'hfd00;
    FD1P3IX pixel_i23 (.D(\Q[8] [23]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[8] [22]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[8] [21]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[8] [20]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[8] [19]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[8] [18]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[8] [17]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[8] [16]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[8] [15]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[8] [14]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[8] [13]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[8] [12]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[8] [11]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[8] [10]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[8] [9]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[8] [8]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[8] [7]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[8] [6]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[8] [5]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[8] [4]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[8] [3]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[8] [2]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[8] [1]), .SP(sclk_c_enable_2418), .CD(n35498), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2385), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2418), 
            .CD(n35498), .CK(sclk_c), .Q(\RdAddress[8] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_2449), .CD(n35469), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_907), .SP(sclk_c_enable_2449), .CD(n35469), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_2449), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=223, LSE_RLINE=223 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 mux_1878_i2_4_lut (.A(n71), .B(n14959[0]), .C(n5853), .D(n52670), 
         .Z(n5854[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i2_4_lut.init = 16'hcfca;
    LUT4 mux_1878_i4_4_lut (.A(n38941), .B(n42484), .C(n5853), .D(n4), 
         .Z(n5854[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut_adj_501 (.A(n42804), .B(n54605), .C(n447[3]), .D(n54723), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut_adj_501.init = 16'hfcee;
    LUT4 mux_1878_i8_4_lut (.A(n5678[7]), .B(n42484), .C(n5853), .D(n54605), 
         .Z(n5854[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i8_4_lut.init = 16'h303a;
    LUT4 mux_1878_i9_4_lut (.A(n5678[8]), .B(n42484), .C(n5853), .D(n54605), 
         .Z(n5854[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i9_4_lut.init = 16'h303a;
    LUT4 mux_1878_i10_4_lut (.A(n80), .B(n42484), .C(n5853), .D(n54605), 
         .Z(n5854[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i10_4_lut.init = 16'h303a;
    LUT4 mux_1878_i13_4_lut (.A(n5678[12]), .B(n42484), .C(n5853), .D(n54605), 
         .Z(n5854[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1878_i13_4_lut.init = 16'h303a;
    PFUMX i38971 (.BLUT(n54995), .ALUT(n54996), .C0(state[1]), .Z(n54997));
    CCU2D add_3118_33 (.A0(bit_counter[31]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48306), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_33.INIT0 = 16'h5999;
    defparam add_3118_33.INIT1 = 16'h0000;
    defparam add_3118_33.INJECT1_0 = "NO";
    defparam add_3118_33.INJECT1_1 = "NO";
    PFUMX i38929 (.BLUT(n54931), .ALUT(n54932), .C0(state[1]), .Z(state_2__N_104[1]));
    CCU2D add_3118_31 (.A0(bit_counter[29]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48305), .COUT(n48306), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_31.INIT0 = 16'h5999;
    defparam add_3118_31.INIT1 = 16'h5999;
    defparam add_3118_31.INJECT1_0 = "NO";
    defparam add_3118_31.INJECT1_1 = "NO";
    CCU2D add_3118_29 (.A0(bit_counter[27]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48304), .COUT(n48305), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_29.INIT0 = 16'h5999;
    defparam add_3118_29.INIT1 = 16'h5999;
    defparam add_3118_29.INJECT1_0 = "NO";
    defparam add_3118_29.INJECT1_1 = "NO";
    CCU2D add_3118_27 (.A0(bit_counter[25]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48303), .COUT(n48304), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_27.INIT0 = 16'h5999;
    defparam add_3118_27.INIT1 = 16'h5999;
    defparam add_3118_27.INJECT1_0 = "NO";
    defparam add_3118_27.INJECT1_1 = "NO";
    CCU2D add_3118_25 (.A0(bit_counter[23]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48302), .COUT(n48303), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_25.INIT0 = 16'h5999;
    defparam add_3118_25.INIT1 = 16'h5999;
    defparam add_3118_25.INJECT1_0 = "NO";
    defparam add_3118_25.INJECT1_1 = "NO";
    CCU2D add_3118_23 (.A0(bit_counter[21]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48301), .COUT(n48302), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_23.INIT0 = 16'h5999;
    defparam add_3118_23.INIT1 = 16'h5999;
    defparam add_3118_23.INJECT1_0 = "NO";
    defparam add_3118_23.INJECT1_1 = "NO";
    CCU2D add_3118_21 (.A0(bit_counter[19]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48300), .COUT(n48301), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_21.INIT0 = 16'h5999;
    defparam add_3118_21.INIT1 = 16'h5999;
    defparam add_3118_21.INJECT1_0 = "NO";
    defparam add_3118_21.INJECT1_1 = "NO";
    CCU2D add_3118_19 (.A0(bit_counter[17]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48299), .COUT(n48300), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_19.INIT0 = 16'h5999;
    defparam add_3118_19.INIT1 = 16'h5999;
    defparam add_3118_19.INJECT1_0 = "NO";
    defparam add_3118_19.INJECT1_1 = "NO";
    CCU2D add_3118_17 (.A0(bit_counter[15]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48298), .COUT(n48299), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_17.INIT0 = 16'h5999;
    defparam add_3118_17.INIT1 = 16'h5999;
    defparam add_3118_17.INJECT1_0 = "NO";
    defparam add_3118_17.INJECT1_1 = "NO";
    CCU2D add_3118_15 (.A0(bit_counter[13]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48297), .COUT(n48298), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_15.INIT0 = 16'h5999;
    defparam add_3118_15.INIT1 = 16'h5999;
    defparam add_3118_15.INJECT1_0 = "NO";
    defparam add_3118_15.INJECT1_1 = "NO";
    CCU2D add_3118_13 (.A0(bit_counter[11]), .B0(n13416), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13416), .C1(GND_net), 
          .D1(GND_net), .CIN(n48296), .COUT(n48297), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3118_13.INIT0 = 16'h5999;
    defparam add_3118_13.INIT1 = 16'h5999;
    defparam add_3118_13.INJECT1_0 = "NO";
    defparam add_3118_13.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module frame_buffer_0
//

module frame_buffer_0 (WrAddress, \RdAddress[9] , Data, \WE[9] , sclk_c, 
            VCC_net, GND_net, \Q[9] ) /* synthesis NGD_DRC_MASK=1 */ ;
    input [8:0]WrAddress;
    input [8:0]\RdAddress[9] ;
    input [23:0]Data;
    input \WE[9] ;
    input sclk_c;
    input VCC_net;
    input GND_net;
    output [23:0]\Q[9] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    PDPW8KC frame_buffer_0_0_1_0 (.DI0(Data[18]), .DI1(Data[19]), .DI2(Data[20]), 
            .DI3(Data[21]), .DI4(Data[22]), .DI5(Data[23]), .DI6(GND_net), 
            .DI7(GND_net), .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), 
            .DI11(GND_net), .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), 
            .DI15(GND_net), .DI16(GND_net), .DI17(GND_net), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[9] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[9] [0]), .ADR5(\RdAddress[9] [1]), 
            .ADR6(\RdAddress[9] [2]), .ADR7(\RdAddress[9] [3]), .ADR8(\RdAddress[9] [4]), 
            .ADR9(\RdAddress[9] [5]), .ADR10(\RdAddress[9] [6]), .ADR11(\RdAddress[9] [7]), 
            .ADR12(\RdAddress[9] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO9(\Q[9] [18]), .DO10(\Q[9] [19]), .DO11(\Q[9] [20]), 
            .DO12(\Q[9] [21]), .DO13(\Q[9] [22]), .DO14(\Q[9] [23])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=229, LSE_RLINE=229 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(229[16:30])
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_1_0.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_1_0.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_1_0.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_1_0.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_1_0.GSR = "ENABLED";
    defparam frame_buffer_0_0_1_0.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_1_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_1_0.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    PDPW8KC frame_buffer_0_0_0_1 (.DI0(Data[0]), .DI1(Data[1]), .DI2(Data[2]), 
            .DI3(Data[3]), .DI4(Data[4]), .DI5(Data[5]), .DI6(Data[6]), 
            .DI7(Data[7]), .DI8(Data[8]), .DI9(Data[9]), .DI10(Data[10]), 
            .DI11(Data[11]), .DI12(Data[12]), .DI13(Data[13]), .DI14(Data[14]), 
            .DI15(Data[15]), .DI16(Data[16]), .DI17(Data[17]), .ADW0(WrAddress[0]), 
            .ADW1(WrAddress[1]), .ADW2(WrAddress[2]), .ADW3(WrAddress[3]), 
            .ADW4(WrAddress[4]), .ADW5(WrAddress[5]), .ADW6(WrAddress[6]), 
            .ADW7(WrAddress[7]), .ADW8(WrAddress[8]), .BE0(VCC_net), .BE1(VCC_net), 
            .CEW(VCC_net), .CLKW(sclk_c), .CSW0(\WE[9] ), .CSW1(GND_net), 
            .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), .ADR2(GND_net), 
            .ADR3(GND_net), .ADR4(\RdAddress[9] [0]), .ADR5(\RdAddress[9] [1]), 
            .ADR6(\RdAddress[9] [2]), .ADR7(\RdAddress[9] [3]), .ADR8(\RdAddress[9] [4]), 
            .ADR9(\RdAddress[9] [5]), .ADR10(\RdAddress[9] [6]), .ADR11(\RdAddress[9] [7]), 
            .ADR12(\RdAddress[9] [8]), .CER(VCC_net), .OCER(VCC_net), 
            .CLKR(sclk_c), .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), 
            .RST(GND_net), .DO0(\Q[9] [9]), .DO1(\Q[9] [10]), .DO2(\Q[9] [11]), 
            .DO3(\Q[9] [12]), .DO4(\Q[9] [13]), .DO5(\Q[9] [14]), .DO6(\Q[9] [15]), 
            .DO7(\Q[9] [16]), .DO8(\Q[9] [17]), .DO9(\Q[9] [0]), .DO10(\Q[9] [1]), 
            .DO11(\Q[9] [2]), .DO12(\Q[9] [3]), .DO13(\Q[9] [4]), .DO14(\Q[9] [5]), 
            .DO15(\Q[9] [6]), .DO16(\Q[9] [7]), .DO17(\Q[9] [8])) /* synthesis MEM_LPC_FILE="frame_buffer_0.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=16, LSE_RCOL=30, LSE_LLINE=229, LSE_RLINE=229 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(229[16:30])
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_W = 18;
    defparam frame_buffer_0_0_0_1.DATA_WIDTH_R = 18;
    defparam frame_buffer_0_0_0_1.REGMODE = "OUTREG";
    defparam frame_buffer_0_0_0_1.CSDECODE_W = "0b001";
    defparam frame_buffer_0_0_0_1.CSDECODE_R = "0b000";
    defparam frame_buffer_0_0_0_1.GSR = "ENABLED";
    defparam frame_buffer_0_0_0_1.RESETMODE = "SYNC";
    defparam frame_buffer_0_0_0_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam frame_buffer_0_0_0_1.INIT_DATA = "STATIC";
    defparam frame_buffer_0_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam frame_buffer_0_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U25 
//

module \WS2812(48000000,"111111111")_U25  (sclk_c, \port_status[3] , ws2813_out_c_3, 
            state, n13101, \Q[3] , \RdAddress[3] , n41629, n10470, 
            GND_net);
    input sclk_c;
    output \port_status[3] ;
    output ws2813_out_c_3;
    output [2:0]state;
    output n13101;
    input [23:0]\Q[3] ;
    output [8:0]\RdAddress[3] ;
    input n41629;
    input n10470;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_889;
    wire [31:0]n7411;
    
    wire sclk_c_enable_35, n54822, sclk_c_enable_36, serial_N_433, sclk_c_enable_39;
    wire [2:0]state_2__N_104;
    
    wire n54956, n42594, n13066, n54955, n53261, n53262;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53263;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1221, n35023;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1209;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1222;
    wire [31:0]bit_counter_31__N_172;
    
    wire n34994, n1, n1_adj_906, n34845;
    wire [31:0]n447;
    
    wire n34841;
    wire [31:0]n7337;
    
    wire n54879, n52974, n52975, n52978, n52976, n52977, n52979, 
        n54616, n54672, n54673, n54729;
    wire [31:0]n7235;
    
    wire serial_N_437;
    wire [6:0]n15022;
    
    wire n42548;
    wire [31:0]bit_counter_31__N_204;
    wire [8:0]n118;
    
    wire n52966, n52967, n15, n14, n52980, n54878, n52973, n54877, 
        n52972, n53260, n53259, n53258, n53257, n52971, n52970, 
        n52969, n52968, n48961, n48960, n48959, n48958, n48957, 
        n48956, n48955, n48954, n48953, n48952, n48951, n48950, 
        n48949, n48948, n48947, n48946, n47613, n47612, n47611, 
        n47610, n47609, n47608, n47607, n47606, n48865, n48864, 
        n48863, n48862, n48861, n48860, n48859, n48858, n48857, 
        n48856, n48855, n48854, n48853, n48852, n48851, n48850, 
        n47605, n47604, n47603, n47602, n48370, n48369, n48368, 
        n48367, n48366, n48365, n48364, n48363, n48362, n48361, 
        n48360, n48359, n48358, n47601, n48357, n48356, n48355, 
        n47600, n47599, n47598, n47596, n47595, n47594, n47593;
    
    FD1P3AX delay_counter_i0_i0 (.D(n7411[0]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54822), .SP(sclk_c_enable_35), .CK(sclk_c), 
            .Q(\port_status[3] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_36), .CK(sclk_c), 
            .Q(ws2813_out_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_39), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_39), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_39), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 mux_2878_i3_then_3_lut (.A(state[2]), .B(state[0]), .C(n13101), 
         .Z(n54956)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam mux_2878_i3_then_3_lut.init = 16'h4040;
    LUT4 mux_2878_i3_else_3_lut (.A(state[2]), .B(state[0]), .C(n42594), 
         .D(n13066), .Z(n54955)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam mux_2878_i3_else_3_lut.init = 16'h4000;
    L6MUX21 i38057 (.D0(n53261), .D1(n53262), .SD(bit_counter[2]), .Z(n53263));
    FD1P3IX pixel_i23 (.D(\Q[3] [23]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[3] [22]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[3] [21]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[3] [20]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[3] [19]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[3] [18]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[3] [17]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[3] [16]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[3] [15]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[3] [14]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[3] [13]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[3] [12]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[3] [11]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[3] [10]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[3] [9]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[3] [8]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[3] [7]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[3] [6]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[3] [5]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[3] [4]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[3] [3]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[3] [2]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[3] [1]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1222), .CD(n34994), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_906), .SP(sclk_c_enable_1222), .CD(n34994), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_889), 
            .CD(n34845), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_889), .CD(n34845), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_889), .CD(n34845), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n7337[4]), .SP(sclk_c_enable_889), .CD(n34841), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54879), .SP(sclk_c_enable_889), .CD(n34841), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    L6MUX21 i37772 (.D0(n52974), .D1(n52975), .SD(bit_counter[2]), .Z(n52978));
    L6MUX21 i37773 (.D0(n52976), .D1(n52977), .SD(bit_counter[2]), .Z(n52979));
    LUT4 i38434_2_lut_rep_801 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1222)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38434_2_lut_rep_801.init = 16'h9999;
    LUT4 i22782_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n34994)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22782_2_lut_2_lut.init = 16'h8888;
    FD1P3AX delay_counter_i0_i1 (.D(n7411[1]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n7411[3]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n7411[7]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n7411[8]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n7411[9]), .SP(sclk_c_enable_889), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n7411[12]), .SP(sclk_c_enable_889), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_613_3_lut (.A(state[2]), .B(n13101), .C(state[1]), 
         .Z(n54616)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_613_3_lut.init = 16'h4040;
    LUT4 i2205_3_lut_rep_669 (.A(state[2]), .B(state[1]), .C(n13101), 
         .Z(n54672)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2205_3_lut_rep_669.init = 16'ha8a8;
    LUT4 i1_2_lut_rep_670 (.A(n13066), .B(n42594), .Z(n54673)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_670.init = 16'h8888;
    LUT4 mux_2177_i1_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[0]), .Z(n7235[0])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_2177_i1_3_lut_4_lut.init = 16'h7f70;
    LUT4 mux_2177_i2_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[1]), .Z(n7235[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_2177_i2_3_lut_4_lut.init = 16'h7f70;
    LUT4 mux_2177_i8_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[7]), .Z(n7235[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_2177_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2177_i9_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[8]), .Z(n7235[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_2177_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2177_i10_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[9]), .Z(n7235[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_2177_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2177_i13_3_lut_4_lut (.A(n13066), .B(n42594), .C(n54729), 
         .D(n447[12]), .Z(n7235[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_2177_i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_1_lut_rep_819 (.A(state[2]), .Z(n54822)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut_rep_819.init = 16'h5555;
    LUT4 i28863_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;
    defparam i28863_3_lut_3_lut.init = 16'h5151;
    LUT4 mux_2193_i1_4_lut (.A(n7235[0]), .B(n15022[0]), .C(n54672), .D(n54616), 
         .Z(n7411[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i1_4_lut.init = 16'hcfca;
    LUT4 i22874_2_lut_2_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n35023)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i22874_2_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i22629_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut (.A(state[1]), .B(n13101), 
         .C(state[2]), .Z(n34841)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i22629_2_lut_3_lut_3_lut_4_lut_3_lut_3_lut.init = 16'he0e0;
    LUT4 i38177_3_lut_rep_716_3_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(sclk_c_enable_1221)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i38177_3_lut_rep_716_3_lut.init = 16'hc1c1;
    LUT4 i38617_2_lut_rep_551_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(n13101), .D(state[2]), .Z(sclk_c_enable_889)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i38617_2_lut_rep_551_2_lut_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13101), .Z(sclk_c_enable_36)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i28688_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15022[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28688_2_lut_3_lut.init = 16'h7070;
    LUT4 i30378_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42548)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i30378_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_726_3_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .Z(n54729)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_726_3_lut.init = 16'h0404;
    LUT4 i37663_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13101), 
         .D(state[1]), .Z(sclk_c_enable_39)) /* synthesis lut_function=(A (C+(D))+!A (B (C+!(D))+!B (C))) */ ;
    defparam i37663_3_lut_4_lut_4_lut_4_lut.init = 16'hfaf4;
    LUT4 i12_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(n13066), 
         .Z(sclk_c_enable_1209)) /* synthesis lut_function=(A (C)+!A !((C+!(D))+!B)) */ ;
    defparam i12_4_lut_4_lut.init = 16'ha4a0;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_417 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_417.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_418 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_418.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_419 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_419.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_420 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_420.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_421 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_421.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_422 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_422.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_423 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_423.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_424 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_424.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_425 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_425.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_426 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_426.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_427 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_427.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_428 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_428.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_429 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_429.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_430 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_430.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_431 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_431.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_432 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_432.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_433 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_433.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_434 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_434.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_435 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_435.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_436 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_436.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_437 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_437.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_438 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_438.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_439 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_439.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_440 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_440.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_441 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_441.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_442 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_442.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_443 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_443.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_444 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_444.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_445 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_445.init = 16'h4040;
    FD1P3IX pixel_i0 (.D(\Q[3] [0]), .SP(sclk_c_enable_1221), .CD(n35023), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1209), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1221), 
            .CD(n35023), .CK(sclk_c), .Q(\RdAddress[3] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1222), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=168, LSE_RLINE=168 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_446 (.A(state[2]), .B(n42594), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_446.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_447 (.A(state[2]), .B(n42594), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_447.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_448 (.A(state[2]), .B(n42594), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_448.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_449 (.A(state[2]), .B(n42594), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_449.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_450 (.A(state[2]), .B(n42594), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_450.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_451 (.A(state[2]), .B(n42594), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_451.init = 16'h1010;
    PFUMX i37768 (.BLUT(n52966), .ALUT(n52967), .C0(bit_counter[1]), .Z(n52974));
    LUT4 i1_2_lut_3_lut_adj_452 (.A(state[2]), .B(n42594), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_452.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_453 (.A(state[2]), .B(n42594), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_453.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_454 (.A(state[2]), .B(n42594), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_454.init = 16'h1010;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[7]), .C(n14), .D(cur_pixel[4]), 
         .Z(n42594)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n52980), .B(n53263), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2878_i1_4_lut (.A(n54673), .B(n41629), .C(n10470), .D(n54729), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2878_i1_4_lut.init = 16'h3a3f;
    LUT4 i6_4_lut (.A(cur_pixel[2]), .B(cur_pixel[8]), .C(cur_pixel[6]), 
         .D(cur_pixel[5]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 mux_2878_i2_4_lut (.A(n13066), .B(n41629), .C(n10470), .D(n54729), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2878_i2_4_lut.init = 16'h3530;
    LUT4 i5_3_lut (.A(cur_pixel[3]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 mux_2183_i3_3_lut_4_lut_then_4_lut (.A(n13101), .B(state[2]), .C(state[0]), 
         .D(n447[2]), .Z(n54878)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (D)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam mux_2183_i3_3_lut_4_lut_then_4_lut.init = 16'hdf02;
    LUT4 i37767_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n52973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37767_3_lut.init = 16'hcaca;
    LUT4 mux_2183_i3_3_lut_4_lut_else_4_lut (.A(state[2]), .B(state[0]), 
         .C(n447[2]), .D(n13066), .Z(n54877)) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam mux_2183_i3_3_lut_4_lut_else_4_lut.init = 16'hb0f4;
    LUT4 i37766_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n52972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37766_3_lut.init = 16'hcaca;
    LUT4 i38054_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38054_3_lut.init = 16'hcaca;
    LUT4 i38053_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38053_3_lut.init = 16'hcaca;
    LUT4 i38052_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38052_3_lut.init = 16'hcaca;
    LUT4 i38051_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38051_3_lut.init = 16'hcaca;
    LUT4 i37765_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n52971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37765_3_lut.init = 16'hcaca;
    LUT4 i37764_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n52970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37764_3_lut.init = 16'hcaca;
    LUT4 i37763_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37763_3_lut.init = 16'hcaca;
    LUT4 i37762_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37762_3_lut.init = 16'hcaca;
    PFUMX i37769 (.BLUT(n52968), .ALUT(n52969), .C0(bit_counter[1]), .Z(n52975));
    LUT4 i37761_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37761_3_lut.init = 16'hcaca;
    PFUMX i37770 (.BLUT(n52970), .ALUT(n52971), .C0(bit_counter[1]), .Z(n52976));
    PFUMX i38055 (.BLUT(n53257), .ALUT(n53258), .C0(bit_counter[1]), .Z(n53261));
    PFUMX i38056 (.BLUT(n53259), .ALUT(n53260), .C0(bit_counter[1]), .Z(n53262));
    LUT4 i28733_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28733_2_lut.init = 16'hbbbb;
    LUT4 i28737_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_906)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28737_2_lut.init = 16'hbbbb;
    PFUMX i37771 (.BLUT(n52972), .ALUT(n52973), .C0(bit_counter[1]), .Z(n52977));
    L6MUX21 i37774 (.D0(n52978), .D1(n52979), .SD(bit_counter[3]), .Z(n52980));
    LUT4 i37760_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37760_3_lut.init = 16'hcaca;
    PFUMX i38893 (.BLUT(n54877), .ALUT(n54878), .C0(state[1]), .Z(n54879));
    LUT4 i22653_4_lut (.A(sclk_c_enable_889), .B(n54616), .C(n54672), 
         .D(n54729), .Z(n34845)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22653_4_lut.init = 16'haaa8;
    LUT4 mux_2183_i5_4_lut (.A(n447[4]), .B(state[0]), .C(n54616), .D(n54729), 
         .Z(n7337[4])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2183_i5_4_lut.init = 16'hc0ca;
    CCU2D add_33929_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48961), 
          .S0(n13101));
    defparam add_33929_cout.INIT0 = 16'h0000;
    defparam add_33929_cout.INIT1 = 16'h0000;
    defparam add_33929_cout.INJECT1_0 = "NO";
    defparam add_33929_cout.INJECT1_1 = "NO";
    CCU2D add_33929_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48960), .COUT(n48961));
    defparam add_33929_31.INIT0 = 16'hf555;
    defparam add_33929_31.INIT1 = 16'h5555;
    defparam add_33929_31.INJECT1_0 = "NO";
    defparam add_33929_31.INJECT1_1 = "NO";
    CCU2D add_33929_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48959), .COUT(n48960));
    defparam add_33929_29.INIT0 = 16'hf555;
    defparam add_33929_29.INIT1 = 16'hf555;
    defparam add_33929_29.INJECT1_0 = "NO";
    defparam add_33929_29.INJECT1_1 = "NO";
    CCU2D add_33929_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48958), .COUT(n48959));
    defparam add_33929_27.INIT0 = 16'hf555;
    defparam add_33929_27.INIT1 = 16'hf555;
    defparam add_33929_27.INJECT1_0 = "NO";
    defparam add_33929_27.INJECT1_1 = "NO";
    CCU2D add_33929_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48957), .COUT(n48958));
    defparam add_33929_25.INIT0 = 16'hf555;
    defparam add_33929_25.INIT1 = 16'hf555;
    defparam add_33929_25.INJECT1_0 = "NO";
    defparam add_33929_25.INJECT1_1 = "NO";
    CCU2D add_33929_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48956), .COUT(n48957));
    defparam add_33929_23.INIT0 = 16'hf555;
    defparam add_33929_23.INIT1 = 16'hf555;
    defparam add_33929_23.INJECT1_0 = "NO";
    defparam add_33929_23.INJECT1_1 = "NO";
    CCU2D add_33929_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48955), .COUT(n48956));
    defparam add_33929_21.INIT0 = 16'hf555;
    defparam add_33929_21.INIT1 = 16'hf555;
    defparam add_33929_21.INJECT1_0 = "NO";
    defparam add_33929_21.INJECT1_1 = "NO";
    CCU2D add_33929_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48954), .COUT(n48955));
    defparam add_33929_19.INIT0 = 16'hf555;
    defparam add_33929_19.INIT1 = 16'hf555;
    defparam add_33929_19.INJECT1_0 = "NO";
    defparam add_33929_19.INJECT1_1 = "NO";
    CCU2D add_33929_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48953), .COUT(n48954));
    defparam add_33929_17.INIT0 = 16'hf555;
    defparam add_33929_17.INIT1 = 16'hf555;
    defparam add_33929_17.INJECT1_0 = "NO";
    defparam add_33929_17.INJECT1_1 = "NO";
    CCU2D add_33929_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48952), .COUT(n48953));
    defparam add_33929_15.INIT0 = 16'hf555;
    defparam add_33929_15.INIT1 = 16'hf555;
    defparam add_33929_15.INJECT1_0 = "NO";
    defparam add_33929_15.INJECT1_1 = "NO";
    CCU2D add_33929_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48951), .COUT(n48952));
    defparam add_33929_13.INIT0 = 16'hf555;
    defparam add_33929_13.INIT1 = 16'hf555;
    defparam add_33929_13.INJECT1_0 = "NO";
    defparam add_33929_13.INJECT1_1 = "NO";
    CCU2D add_33929_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48950), .COUT(n48951));
    defparam add_33929_11.INIT0 = 16'hf555;
    defparam add_33929_11.INIT1 = 16'hf555;
    defparam add_33929_11.INJECT1_0 = "NO";
    defparam add_33929_11.INJECT1_1 = "NO";
    CCU2D add_33929_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48949), .COUT(n48950));
    defparam add_33929_9.INIT0 = 16'hf555;
    defparam add_33929_9.INIT1 = 16'hf555;
    defparam add_33929_9.INJECT1_0 = "NO";
    defparam add_33929_9.INJECT1_1 = "NO";
    CCU2D add_33929_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48948), .COUT(n48949));
    defparam add_33929_7.INIT0 = 16'hf555;
    defparam add_33929_7.INIT1 = 16'hf555;
    defparam add_33929_7.INJECT1_0 = "NO";
    defparam add_33929_7.INJECT1_1 = "NO";
    CCU2D add_33929_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48947), .COUT(n48948));
    defparam add_33929_5.INIT0 = 16'hf555;
    defparam add_33929_5.INIT1 = 16'hf555;
    defparam add_33929_5.INJECT1_0 = "NO";
    defparam add_33929_5.INJECT1_1 = "NO";
    CCU2D add_33929_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48946), .COUT(n48947));
    defparam add_33929_3.INIT0 = 16'hf555;
    defparam add_33929_3.INIT1 = 16'hf555;
    defparam add_33929_3.INJECT1_0 = "NO";
    defparam add_33929_3.INJECT1_1 = "NO";
    CCU2D add_33929_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48946));
    defparam add_33929_1.INIT0 = 16'hF000;
    defparam add_33929_1.INIT1 = 16'ha666;
    defparam add_33929_1.INJECT1_0 = "NO";
    defparam add_33929_1.INJECT1_1 = "NO";
    LUT4 mux_2193_i2_4_lut (.A(n7235[1]), .B(n15022[0]), .C(n54672), .D(n54616), 
         .Z(n7411[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2193_i4_4_lut (.A(n7235[3]), .B(n42548), .C(n54672), .D(n54616), 
         .Z(n7411[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i4_4_lut.init = 16'h3f3a;
    LUT4 mux_2177_i4_4_lut (.A(n447[3]), .B(n42594), .C(n54729), .D(n13066), 
         .Z(n7235[3])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2177_i4_4_lut.init = 16'hcafa;
    LUT4 mux_2193_i8_4_lut (.A(n7235[7]), .B(n42548), .C(n54672), .D(n54616), 
         .Z(n7411[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i8_4_lut.init = 16'h303a;
    LUT4 mux_2193_i9_4_lut (.A(n7235[8]), .B(n42548), .C(n54672), .D(n54616), 
         .Z(n7411[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i9_4_lut.init = 16'h303a;
    LUT4 mux_2193_i10_4_lut (.A(n7235[9]), .B(n42548), .C(n54672), .D(n54616), 
         .Z(n7411[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i10_4_lut.init = 16'h303a;
    LUT4 mux_2193_i13_4_lut (.A(n7235[12]), .B(n42548), .C(n54672), .D(n54616), 
         .Z(n7411[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2193_i13_4_lut.init = 16'h303a;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47613), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47612), .COUT(n47613), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47611), .COUT(n47612), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47610), .COUT(n47611), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47609), .COUT(n47610), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47608), .COUT(n47609), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47607), .COUT(n47608), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47606), .COUT(n47607), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_33934_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48865), 
          .S0(n13066));
    defparam add_33934_cout.INIT0 = 16'h0000;
    defparam add_33934_cout.INIT1 = 16'h0000;
    defparam add_33934_cout.INJECT1_0 = "NO";
    defparam add_33934_cout.INJECT1_1 = "NO";
    CCU2D add_33934_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48864), .COUT(n48865));
    defparam add_33934_31.INIT0 = 16'hf555;
    defparam add_33934_31.INIT1 = 16'h5555;
    defparam add_33934_31.INJECT1_0 = "NO";
    defparam add_33934_31.INJECT1_1 = "NO";
    CCU2D add_33934_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48863), .COUT(n48864));
    defparam add_33934_29.INIT0 = 16'hf555;
    defparam add_33934_29.INIT1 = 16'hf555;
    defparam add_33934_29.INJECT1_0 = "NO";
    defparam add_33934_29.INJECT1_1 = "NO";
    CCU2D add_33934_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48862), .COUT(n48863));
    defparam add_33934_27.INIT0 = 16'hf555;
    defparam add_33934_27.INIT1 = 16'hf555;
    defparam add_33934_27.INJECT1_0 = "NO";
    defparam add_33934_27.INJECT1_1 = "NO";
    CCU2D add_33934_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48861), .COUT(n48862));
    defparam add_33934_25.INIT0 = 16'hf555;
    defparam add_33934_25.INIT1 = 16'hf555;
    defparam add_33934_25.INJECT1_0 = "NO";
    defparam add_33934_25.INJECT1_1 = "NO";
    CCU2D add_33934_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48860), .COUT(n48861));
    defparam add_33934_23.INIT0 = 16'hf555;
    defparam add_33934_23.INIT1 = 16'hf555;
    defparam add_33934_23.INJECT1_0 = "NO";
    defparam add_33934_23.INJECT1_1 = "NO";
    CCU2D add_33934_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48859), .COUT(n48860));
    defparam add_33934_21.INIT0 = 16'hf555;
    defparam add_33934_21.INIT1 = 16'hf555;
    defparam add_33934_21.INJECT1_0 = "NO";
    defparam add_33934_21.INJECT1_1 = "NO";
    CCU2D add_33934_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48858), .COUT(n48859));
    defparam add_33934_19.INIT0 = 16'hf555;
    defparam add_33934_19.INIT1 = 16'hf555;
    defparam add_33934_19.INJECT1_0 = "NO";
    defparam add_33934_19.INJECT1_1 = "NO";
    CCU2D add_33934_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48857), .COUT(n48858));
    defparam add_33934_17.INIT0 = 16'hf555;
    defparam add_33934_17.INIT1 = 16'hf555;
    defparam add_33934_17.INJECT1_0 = "NO";
    defparam add_33934_17.INJECT1_1 = "NO";
    CCU2D add_33934_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48856), .COUT(n48857));
    defparam add_33934_15.INIT0 = 16'hf555;
    defparam add_33934_15.INIT1 = 16'hf555;
    defparam add_33934_15.INJECT1_0 = "NO";
    defparam add_33934_15.INJECT1_1 = "NO";
    CCU2D add_33934_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48855), .COUT(n48856));
    defparam add_33934_13.INIT0 = 16'hf555;
    defparam add_33934_13.INIT1 = 16'hf555;
    defparam add_33934_13.INJECT1_0 = "NO";
    defparam add_33934_13.INJECT1_1 = "NO";
    CCU2D add_33934_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48854), .COUT(n48855));
    defparam add_33934_11.INIT0 = 16'hf555;
    defparam add_33934_11.INIT1 = 16'hf555;
    defparam add_33934_11.INJECT1_0 = "NO";
    defparam add_33934_11.INJECT1_1 = "NO";
    CCU2D add_33934_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48853), .COUT(n48854));
    defparam add_33934_9.INIT0 = 16'hf555;
    defparam add_33934_9.INIT1 = 16'hf555;
    defparam add_33934_9.INJECT1_0 = "NO";
    defparam add_33934_9.INJECT1_1 = "NO";
    CCU2D add_33934_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48852), .COUT(n48853));
    defparam add_33934_7.INIT0 = 16'hf555;
    defparam add_33934_7.INIT1 = 16'hf555;
    defparam add_33934_7.INJECT1_0 = "NO";
    defparam add_33934_7.INJECT1_1 = "NO";
    CCU2D add_33934_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48851), .COUT(n48852));
    defparam add_33934_5.INIT0 = 16'hf555;
    defparam add_33934_5.INIT1 = 16'hf555;
    defparam add_33934_5.INJECT1_0 = "NO";
    defparam add_33934_5.INJECT1_1 = "NO";
    CCU2D add_33934_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48850), .COUT(n48851));
    defparam add_33934_3.INIT0 = 16'hf555;
    defparam add_33934_3.INIT1 = 16'hf555;
    defparam add_33934_3.INJECT1_0 = "NO";
    defparam add_33934_3.INJECT1_1 = "NO";
    CCU2D add_33934_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48850));
    defparam add_33934_1.INIT0 = 16'hF000;
    defparam add_33934_1.INIT1 = 16'ha666;
    defparam add_33934_1.INJECT1_0 = "NO";
    defparam add_33934_1.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47605), .COUT(n47606), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47604), .COUT(n47605), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47603), .COUT(n47604), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47602), .COUT(n47603), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_3108_33 (.A0(bit_counter[31]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48370), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_33.INIT0 = 16'h5999;
    defparam add_3108_33.INIT1 = 16'h0000;
    defparam add_3108_33.INJECT1_0 = "NO";
    defparam add_3108_33.INJECT1_1 = "NO";
    CCU2D add_3108_31 (.A0(bit_counter[29]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48369), .COUT(n48370), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_31.INIT0 = 16'h5999;
    defparam add_3108_31.INIT1 = 16'h5999;
    defparam add_3108_31.INJECT1_0 = "NO";
    defparam add_3108_31.INJECT1_1 = "NO";
    CCU2D add_3108_29 (.A0(bit_counter[27]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48368), .COUT(n48369), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_29.INIT0 = 16'h5999;
    defparam add_3108_29.INIT1 = 16'h5999;
    defparam add_3108_29.INJECT1_0 = "NO";
    defparam add_3108_29.INJECT1_1 = "NO";
    CCU2D add_3108_27 (.A0(bit_counter[25]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48367), .COUT(n48368), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_27.INIT0 = 16'h5999;
    defparam add_3108_27.INIT1 = 16'h5999;
    defparam add_3108_27.INJECT1_0 = "NO";
    defparam add_3108_27.INJECT1_1 = "NO";
    CCU2D add_3108_25 (.A0(bit_counter[23]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48366), .COUT(n48367), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_25.INIT0 = 16'h5999;
    defparam add_3108_25.INIT1 = 16'h5999;
    defparam add_3108_25.INJECT1_0 = "NO";
    defparam add_3108_25.INJECT1_1 = "NO";
    CCU2D add_3108_23 (.A0(bit_counter[21]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48365), .COUT(n48366), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_23.INIT0 = 16'h5999;
    defparam add_3108_23.INIT1 = 16'h5999;
    defparam add_3108_23.INJECT1_0 = "NO";
    defparam add_3108_23.INJECT1_1 = "NO";
    CCU2D add_3108_21 (.A0(bit_counter[19]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48364), .COUT(n48365), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_21.INIT0 = 16'h5999;
    defparam add_3108_21.INIT1 = 16'h5999;
    defparam add_3108_21.INJECT1_0 = "NO";
    defparam add_3108_21.INJECT1_1 = "NO";
    CCU2D add_3108_19 (.A0(bit_counter[17]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48363), .COUT(n48364), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_19.INIT0 = 16'h5999;
    defparam add_3108_19.INIT1 = 16'h5999;
    defparam add_3108_19.INJECT1_0 = "NO";
    defparam add_3108_19.INJECT1_1 = "NO";
    CCU2D add_3108_17 (.A0(bit_counter[15]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48362), .COUT(n48363), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_17.INIT0 = 16'h5999;
    defparam add_3108_17.INIT1 = 16'h5999;
    defparam add_3108_17.INJECT1_0 = "NO";
    defparam add_3108_17.INJECT1_1 = "NO";
    CCU2D add_3108_15 (.A0(bit_counter[13]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48361), .COUT(n48362), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_15.INIT0 = 16'h5999;
    defparam add_3108_15.INIT1 = 16'h5999;
    defparam add_3108_15.INJECT1_0 = "NO";
    defparam add_3108_15.INJECT1_1 = "NO";
    CCU2D add_3108_13 (.A0(bit_counter[11]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48360), .COUT(n48361), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_13.INIT0 = 16'h5999;
    defparam add_3108_13.INIT1 = 16'h5999;
    defparam add_3108_13.INJECT1_0 = "NO";
    defparam add_3108_13.INJECT1_1 = "NO";
    CCU2D add_3108_11 (.A0(bit_counter[9]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48359), .COUT(n48360), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_11.INIT0 = 16'h5999;
    defparam add_3108_11.INIT1 = 16'h5999;
    defparam add_3108_11.INJECT1_0 = "NO";
    defparam add_3108_11.INJECT1_1 = "NO";
    CCU2D add_3108_9 (.A0(bit_counter[7]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48358), .COUT(n48359), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_9.INIT0 = 16'h5999;
    defparam add_3108_9.INIT1 = 16'h5999;
    defparam add_3108_9.INJECT1_0 = "NO";
    defparam add_3108_9.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47601), .COUT(n47602), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_3108_7 (.A0(bit_counter[5]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48357), .COUT(n48358), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_7.INIT0 = 16'h5999;
    defparam add_3108_7.INIT1 = 16'h5999;
    defparam add_3108_7.INJECT1_0 = "NO";
    defparam add_3108_7.INJECT1_1 = "NO";
    CCU2D add_3108_5 (.A0(bit_counter[3]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48356), .COUT(n48357), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_5.INIT0 = 16'h5999;
    defparam add_3108_5.INIT1 = 16'h5999;
    defparam add_3108_5.INJECT1_0 = "NO";
    defparam add_3108_5.INJECT1_1 = "NO";
    CCU2D add_3108_3 (.A0(bit_counter[1]), .B0(n13066), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13066), .C1(GND_net), 
          .D1(GND_net), .CIN(n48355), .COUT(n48356), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_3.INIT0 = 16'h5999;
    defparam add_3108_3.INIT1 = 16'h5999;
    defparam add_3108_3.INJECT1_0 = "NO";
    defparam add_3108_3.INJECT1_1 = "NO";
    CCU2D add_3108_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13066), .C1(GND_net), .D1(GND_net), 
          .COUT(n48355), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3108_1.INIT0 = 16'hF000;
    defparam add_3108_1.INIT1 = 16'h5999;
    defparam add_3108_1.INJECT1_0 = "NO";
    defparam add_3108_1.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47600), .COUT(n47601), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47599), .COUT(n47600), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47598), .COUT(n47599), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47598), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47596), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47595), .COUT(n47596), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47594), .COUT(n47595), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47593), .COUT(n47594), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47593), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    PFUMX i38945 (.BLUT(n54955), .ALUT(n54956), .C0(state[1]), .Z(state_2__N_104[2]));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U22 
//

module \WS2812(48000000,"111111111")_U22  (sclk_c, \port_status[6] , ws2813_out_c_6, 
            \Q[6] , \RdAddress[6] , GND_net);
    input sclk_c;
    output \port_status[6] ;
    output ws2813_out_c_6;
    input [23:0]\Q[6] ;
    output [8:0]\RdAddress[6] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n53019, n53020;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53023, n53021, n53022, n53024;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_939;
    wire [31:0]n6076;
    
    wire sclk_c_enable_61, n54811, sclk_c_enable_62, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_66;
    wire [2:0]state_2__N_104;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1185, n35308;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1184;
    wire [8:0]cur_pixel_8__N_107;
    
    wire n13311, sclk_c_enable_1186;
    wire [31:0]bit_counter_31__N_172;
    
    wire n9669, n35279, n1, n1_adj_905;
    wire [31:0]n447;
    
    wire n54926, n54925, n54941, n13276, n54940, n53282, n53283, 
        n53284, n35130, n35126, n54927, n54942, n54666, n54612, 
        n42584, n54667, n54604, n54726, n103, serial_N_437, n54821;
    wire [31:0]n5900;
    
    wire n76, n54722;
    wire [6:0]n14767;
    
    wire n69, n68, n39205;
    wire [31:0]bit_counter_31__N_204;
    
    wire n53011, n53012, n53013, n53014, n53015, n53016, n53017, 
        n53018, n6075, n52721;
    wire [8:0]n118;
    
    wire n15, n14, n53025, n53281, n53280, n53279, n53278, n48529, 
        n48528, n48527, n48526, n48525, n48524, n48523, n48522, 
        n48521, n48520, n48519, n48518, n48517, n48516, n48515, 
        n48514, n4, n47708, n47707, n47706, n47705, n47704, n47703, 
        n47702, n47701, n47700, n48801, n48800, n48799, n48798, 
        n48797, n48796, n48795, n48794, n48793, n48792, n48791, 
        n48790, n48789, n48788, n48787, n48786, n47699, n47698, 
        n47697, n47696, n47695, n47694, n47693, n47691, n47690, 
        n48322, n47689, n47688, n48321, n48320, n48319, n48318, 
        n48317, n48316, n48315, n48314, n48313, n48312, n48311, 
        n48310, n48309, n48308, n48307;
    
    L6MUX21 i37817 (.D0(n53019), .D1(n53020), .SD(bit_counter[2]), .Z(n53023));
    L6MUX21 i37818 (.D0(n53021), .D1(n53022), .SD(bit_counter[2]), .Z(n53024));
    FD1P3AX delay_counter_i0_i0 (.D(n6076[0]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54811), .SP(sclk_c_enable_61), .CK(sclk_c), 
            .Q(\port_status[6] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_62), .CK(sclk_c), 
            .Q(ws2813_out_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_66), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_66), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_66), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    FD1P3IX pixel_i23 (.D(\Q[6] [23]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[6] [22]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[6] [21]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[6] [20]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[6] [19]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[6] [18]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[6] [17]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[6] [16]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[6] [15]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[6] [14]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[6] [13]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[6] [12]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[6] [11]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[6] [10]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[6] [9]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[6] [8]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[6] [7]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[6] [6]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[6] [5]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[6] [4]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[6] [3]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[6] [2]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[6] [1]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    LUT4 i38453_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13311), .Z(sclk_c_enable_66)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38453_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13311), .Z(n9669)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1186), .CD(n35279), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_905), .SP(sclk_c_enable_1186), .CD(n35279), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 mux_1898_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13311), .Z(n54926)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_1898_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_1898_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13311), .Z(n54925)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_1898_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 mux_1898_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13311), .Z(n54941)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1898_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_1898_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13276), .Z(n54940)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1898_i3_4_lut_else_4_lut.init = 16'hd0f2;
    L6MUX21 i38078 (.D0(n53282), .D1(n53283), .SD(bit_counter[2]), .Z(n53284));
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_939), 
            .CD(n35130), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_939), .CD(n35130), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_939), .CD(n35130), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54927), .SP(sclk_c_enable_939), .CD(n35126), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54942), .SP(sclk_c_enable_939), .CD(n35126), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_663 (.A(state[2]), .B(n13311), .Z(n54666)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_663.init = 16'h4444;
    LUT4 i1_2_lut_rep_609_3_lut (.A(state[2]), .B(n13311), .C(state[1]), 
         .Z(n54612)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_609_3_lut.init = 16'h4040;
    LUT4 i38610_3_lut_rep_610_4_lut (.A(state[2]), .B(n13311), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_939)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38610_3_lut_rep_610_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_rep_664 (.A(n42584), .B(n13276), .Z(n54667)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_664.init = 16'h8888;
    LUT4 i1_2_lut_rep_601_3_lut (.A(n42584), .B(n13276), .C(state[1]), 
         .Z(n54604)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_601_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42584), .B(n13276), .C(n54726), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 i27012_1_lut_rep_808 (.A(state[2]), .Z(n54811)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27012_1_lut_rep_808.init = 16'h5555;
    LUT4 i28914_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28914_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_3_lut_4_lut (.A(n54604), .B(n54821), .C(n447[7]), .D(n54726), 
         .Z(n5900[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_374 (.A(n54604), .B(n54821), .C(n447[8]), 
         .D(n54726), .Z(n5900[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_374.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_375 (.A(n54604), .B(n54821), .C(n447[9]), 
         .D(n54726), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_375.init = 16'hf888;
    FD1P3AX delay_counter_i0_i1 (.D(n6076[1]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n6076[3]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n6076[7]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n6076[8]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n6076[9]), .SP(sclk_c_enable_939), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n6076[12]), .SP(sclk_c_enable_939), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_719_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54722)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_719_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n14767[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_723_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54726)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_723_3_lut.init = 16'hefef;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n13311), 
         .Z(sclk_c_enable_62)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_3_lut_rep_699_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_1185)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_699_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_376 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_376.init = 16'he0f0;
    LUT4 i23159_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n35308)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i23159_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_818 (.A(state[2]), .B(state[0]), .Z(n54821)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_818.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_377 (.A(state[2]), .B(state[0]), .C(n13276), 
         .D(state[1]), .Z(n39205)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_377.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n13276), 
         .D(state[1]), .Z(sclk_c_enable_1184)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_3_lut_adj_378 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_378.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_379 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_379.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_380 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_380.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_381 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_381.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_382 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_382.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_383 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_383.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_384 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_384.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_385 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_385.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_386 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_386.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_387 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_387.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_388 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_388.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_389 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_389.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_390 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_390.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_391 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_391.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_392 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_392.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_393 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_393.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_394 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_394.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_395 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_395.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_396 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_396.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_397 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_397.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_398 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_398.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_399 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_399.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_400 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_400.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_401 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_401.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_402 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_402.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_403 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_403.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_404 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_404.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_405 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_405.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_406 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_406.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_407 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_407.init = 16'h4040;
    PFUMX i37813 (.BLUT(n53011), .ALUT(n53012), .C0(bit_counter[1]), .Z(n53019));
    PFUMX i37814 (.BLUT(n53013), .ALUT(n53014), .C0(bit_counter[1]), .Z(n53020));
    LUT4 i38410_2_lut_rep_826 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1186)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38410_2_lut_rep_826.init = 16'h9999;
    LUT4 i23067_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35279)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23067_2_lut_2_lut.init = 16'h8888;
    PFUMX i37815 (.BLUT(n53015), .ALUT(n53016), .C0(bit_counter[1]), .Z(n53021));
    LUT4 i28768_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28768_2_lut.init = 16'hbbbb;
    LUT4 i28767_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_905)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28767_2_lut.init = 16'hbbbb;
    FD1P3IX pixel_i0 (.D(\Q[6] [0]), .SP(sclk_c_enable_1185), .CD(n35308), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1184), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1185), 
            .CD(n35308), .CK(sclk_c), .Q(\RdAddress[6] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1186), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=201, LSE_RLINE=201 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    PFUMX i37816 (.BLUT(n53017), .ALUT(n53018), .C0(bit_counter[1]), .Z(n53022));
    LUT4 mux_2707_i2_4_lut_4_lut (.A(n54722), .B(n54726), .C(n9669), .D(n13276), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2707_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 mux_1908_i1_4_lut (.A(n69), .B(n14767[0]), .C(n6075), .D(n52721), 
         .Z(n6076[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i1_4_lut.init = 16'hcfca;
    LUT4 i1_2_lut_3_lut_adj_408 (.A(state[2]), .B(n42584), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_408.init = 16'h1010;
    LUT4 i1920_3_lut (.A(state[2]), .B(state[1]), .C(n13311), .Z(n6075)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1920_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_3_lut_adj_409 (.A(state[2]), .B(n42584), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_409.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_410 (.A(state[2]), .B(n42584), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_410.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_411 (.A(state[2]), .B(n42584), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_411.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_412 (.A(state[2]), .B(n42584), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_412.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_413 (.A(state[2]), .B(n42584), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_413.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_414 (.A(state[2]), .B(n42584), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_414.init = 16'h1010;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[2]), .C(n14), .D(cur_pixel[8]), 
         .Z(n42584)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[3]), .B(cur_pixel[5]), .C(cur_pixel[7]), 
         .D(cur_pixel[4]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[6]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_415 (.A(state[2]), .B(n42584), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_415.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_416 (.A(state[2]), .B(n42584), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_416.init = 16'h1010;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53025), .B(n53284), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2707_i1_4_lut (.A(n54667), .B(n54722), .C(n9669), .D(n54726), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2707_i1_4_lut.init = 16'h3f3a;
    LUT4 i38075_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38075_3_lut.init = 16'hcaca;
    LUT4 i38074_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38074_3_lut.init = 16'hcaca;
    LUT4 i38073_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38073_3_lut.init = 16'hcaca;
    LUT4 i38072_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38072_3_lut.init = 16'hcaca;
    LUT4 i22938_4_lut (.A(sclk_c_enable_939), .B(n54726), .C(n6075), .D(n54612), 
         .Z(n35130)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22938_4_lut.init = 16'haaa2;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54821), .B(state[1]), .C(n54667), .D(n54666), 
         .Z(n52721)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    L6MUX21 i37819 (.D0(n53023), .D1(n53024), .SD(bit_counter[3]), .Z(n53025));
    CCU2D add_33898_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48529), 
          .S0(n13311));
    defparam add_33898_cout.INIT0 = 16'h0000;
    defparam add_33898_cout.INIT1 = 16'h0000;
    defparam add_33898_cout.INJECT1_0 = "NO";
    defparam add_33898_cout.INJECT1_1 = "NO";
    CCU2D add_33898_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48528), .COUT(n48529));
    defparam add_33898_31.INIT0 = 16'hf555;
    defparam add_33898_31.INIT1 = 16'h5555;
    defparam add_33898_31.INJECT1_0 = "NO";
    defparam add_33898_31.INJECT1_1 = "NO";
    CCU2D add_33898_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48527), .COUT(n48528));
    defparam add_33898_29.INIT0 = 16'hf555;
    defparam add_33898_29.INIT1 = 16'hf555;
    defparam add_33898_29.INJECT1_0 = "NO";
    defparam add_33898_29.INJECT1_1 = "NO";
    CCU2D add_33898_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48526), .COUT(n48527));
    defparam add_33898_27.INIT0 = 16'hf555;
    defparam add_33898_27.INIT1 = 16'hf555;
    defparam add_33898_27.INJECT1_0 = "NO";
    defparam add_33898_27.INJECT1_1 = "NO";
    CCU2D add_33898_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48525), .COUT(n48526));
    defparam add_33898_25.INIT0 = 16'hf555;
    defparam add_33898_25.INIT1 = 16'hf555;
    defparam add_33898_25.INJECT1_0 = "NO";
    defparam add_33898_25.INJECT1_1 = "NO";
    CCU2D add_33898_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48524), .COUT(n48525));
    defparam add_33898_23.INIT0 = 16'hf555;
    defparam add_33898_23.INIT1 = 16'hf555;
    defparam add_33898_23.INJECT1_0 = "NO";
    defparam add_33898_23.INJECT1_1 = "NO";
    CCU2D add_33898_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48523), .COUT(n48524));
    defparam add_33898_21.INIT0 = 16'hf555;
    defparam add_33898_21.INIT1 = 16'hf555;
    defparam add_33898_21.INJECT1_0 = "NO";
    defparam add_33898_21.INJECT1_1 = "NO";
    CCU2D add_33898_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48522), .COUT(n48523));
    defparam add_33898_19.INIT0 = 16'hf555;
    defparam add_33898_19.INIT1 = 16'hf555;
    defparam add_33898_19.INJECT1_0 = "NO";
    defparam add_33898_19.INJECT1_1 = "NO";
    CCU2D add_33898_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48521), .COUT(n48522));
    defparam add_33898_17.INIT0 = 16'hf555;
    defparam add_33898_17.INIT1 = 16'hf555;
    defparam add_33898_17.INJECT1_0 = "NO";
    defparam add_33898_17.INJECT1_1 = "NO";
    CCU2D add_33898_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48520), .COUT(n48521));
    defparam add_33898_15.INIT0 = 16'hf555;
    defparam add_33898_15.INIT1 = 16'hf555;
    defparam add_33898_15.INJECT1_0 = "NO";
    defparam add_33898_15.INJECT1_1 = "NO";
    PFUMX i38076 (.BLUT(n53278), .ALUT(n53279), .C0(bit_counter[1]), .Z(n53282));
    PFUMX i38077 (.BLUT(n53280), .ALUT(n53281), .C0(bit_counter[1]), .Z(n53283));
    CCU2D add_33898_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48519), .COUT(n48520));
    defparam add_33898_13.INIT0 = 16'hf555;
    defparam add_33898_13.INIT1 = 16'hf555;
    defparam add_33898_13.INJECT1_0 = "NO";
    defparam add_33898_13.INJECT1_1 = "NO";
    CCU2D add_33898_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48518), .COUT(n48519));
    defparam add_33898_11.INIT0 = 16'hf555;
    defparam add_33898_11.INIT1 = 16'hf555;
    defparam add_33898_11.INJECT1_0 = "NO";
    defparam add_33898_11.INJECT1_1 = "NO";
    CCU2D add_33898_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48517), .COUT(n48518));
    defparam add_33898_9.INIT0 = 16'hf555;
    defparam add_33898_9.INIT1 = 16'hf555;
    defparam add_33898_9.INJECT1_0 = "NO";
    defparam add_33898_9.INJECT1_1 = "NO";
    CCU2D add_33898_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48516), .COUT(n48517));
    defparam add_33898_7.INIT0 = 16'hf555;
    defparam add_33898_7.INIT1 = 16'hf555;
    defparam add_33898_7.INJECT1_0 = "NO";
    defparam add_33898_7.INJECT1_1 = "NO";
    CCU2D add_33898_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48515), .COUT(n48516));
    defparam add_33898_5.INIT0 = 16'hf555;
    defparam add_33898_5.INIT1 = 16'hf555;
    defparam add_33898_5.INJECT1_0 = "NO";
    defparam add_33898_5.INJECT1_1 = "NO";
    CCU2D add_33898_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48514), .COUT(n48515));
    defparam add_33898_3.INIT0 = 16'hf555;
    defparam add_33898_3.INIT1 = 16'hf555;
    defparam add_33898_3.INJECT1_0 = "NO";
    defparam add_33898_3.INJECT1_1 = "NO";
    CCU2D add_33898_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48514));
    defparam add_33898_1.INIT0 = 16'hF000;
    defparam add_33898_1.INIT1 = 16'ha666;
    defparam add_33898_1.INJECT1_0 = "NO";
    defparam add_33898_1.INJECT1_1 = "NO";
    LUT4 i37812_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37812_3_lut.init = 16'hcaca;
    LUT4 i37811_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37811_3_lut.init = 16'hcaca;
    LUT4 i37810_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37810_3_lut.init = 16'hcaca;
    LUT4 i37809_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37809_3_lut.init = 16'hcaca;
    LUT4 i37808_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37808_3_lut.init = 16'hcaca;
    LUT4 i37807_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37807_3_lut.init = 16'hcaca;
    LUT4 i37806_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37806_3_lut.init = 16'hcaca;
    LUT4 i37805_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37805_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54667), .C(n13311), .D(n54821), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    LUT4 mux_1908_i2_4_lut (.A(n68), .B(n14767[0]), .C(n6075), .D(n52721), 
         .Z(n6076[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i2_4_lut.init = 16'hcfca;
    LUT4 mux_1908_i4_4_lut (.A(n39205), .B(n54722), .C(n6075), .D(n4), 
         .Z(n6076[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42584), .B(n54612), .C(n447[3]), .D(n54726), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_1908_i8_4_lut (.A(n5900[7]), .B(n54722), .C(n6075), .D(n54612), 
         .Z(n6076[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i8_4_lut.init = 16'h303a;
    LUT4 i22914_2_lut_4_lut (.A(n54666), .B(state[0]), .C(state[1]), .D(n6075), 
         .Z(n35126)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i22914_2_lut_4_lut.init = 16'hfd00;
    LUT4 mux_1908_i9_4_lut (.A(n5900[8]), .B(n54722), .C(n6075), .D(n54612), 
         .Z(n6076[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i9_4_lut.init = 16'h303a;
    LUT4 mux_1908_i10_4_lut (.A(n76), .B(n54722), .C(n6075), .D(n54612), 
         .Z(n6076[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i10_4_lut.init = 16'h303a;
    LUT4 mux_1908_i13_4_lut (.A(n54612), .B(n54722), .C(n6075), .D(n103), 
         .Z(n6076[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1908_i13_4_lut.init = 16'h3530;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47708), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47707), .COUT(n47708), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47706), .COUT(n47707), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47705), .COUT(n47706), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47704), .COUT(n47705), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47703), .COUT(n47704), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47702), .COUT(n47703), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47701), .COUT(n47702), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47700), .COUT(n47701), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_33905_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48801), 
          .S0(n13276));
    defparam add_33905_cout.INIT0 = 16'h0000;
    defparam add_33905_cout.INIT1 = 16'h0000;
    defparam add_33905_cout.INJECT1_0 = "NO";
    defparam add_33905_cout.INJECT1_1 = "NO";
    CCU2D add_33905_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48800), .COUT(n48801));
    defparam add_33905_31.INIT0 = 16'hf555;
    defparam add_33905_31.INIT1 = 16'h5555;
    defparam add_33905_31.INJECT1_0 = "NO";
    defparam add_33905_31.INJECT1_1 = "NO";
    CCU2D add_33905_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48799), .COUT(n48800));
    defparam add_33905_29.INIT0 = 16'hf555;
    defparam add_33905_29.INIT1 = 16'hf555;
    defparam add_33905_29.INJECT1_0 = "NO";
    defparam add_33905_29.INJECT1_1 = "NO";
    CCU2D add_33905_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48798), .COUT(n48799));
    defparam add_33905_27.INIT0 = 16'hf555;
    defparam add_33905_27.INIT1 = 16'hf555;
    defparam add_33905_27.INJECT1_0 = "NO";
    defparam add_33905_27.INJECT1_1 = "NO";
    CCU2D add_33905_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48797), .COUT(n48798));
    defparam add_33905_25.INIT0 = 16'hf555;
    defparam add_33905_25.INIT1 = 16'hf555;
    defparam add_33905_25.INJECT1_0 = "NO";
    defparam add_33905_25.INJECT1_1 = "NO";
    CCU2D add_33905_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48796), .COUT(n48797));
    defparam add_33905_23.INIT0 = 16'hf555;
    defparam add_33905_23.INIT1 = 16'hf555;
    defparam add_33905_23.INJECT1_0 = "NO";
    defparam add_33905_23.INJECT1_1 = "NO";
    CCU2D add_33905_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48795), .COUT(n48796));
    defparam add_33905_21.INIT0 = 16'hf555;
    defparam add_33905_21.INIT1 = 16'hf555;
    defparam add_33905_21.INJECT1_0 = "NO";
    defparam add_33905_21.INJECT1_1 = "NO";
    CCU2D add_33905_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48794), .COUT(n48795));
    defparam add_33905_19.INIT0 = 16'hf555;
    defparam add_33905_19.INIT1 = 16'hf555;
    defparam add_33905_19.INJECT1_0 = "NO";
    defparam add_33905_19.INJECT1_1 = "NO";
    CCU2D add_33905_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48793), .COUT(n48794));
    defparam add_33905_17.INIT0 = 16'hf555;
    defparam add_33905_17.INIT1 = 16'hf555;
    defparam add_33905_17.INJECT1_0 = "NO";
    defparam add_33905_17.INJECT1_1 = "NO";
    CCU2D add_33905_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48792), .COUT(n48793));
    defparam add_33905_15.INIT0 = 16'hf555;
    defparam add_33905_15.INIT1 = 16'hf555;
    defparam add_33905_15.INJECT1_0 = "NO";
    defparam add_33905_15.INJECT1_1 = "NO";
    CCU2D add_33905_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48791), .COUT(n48792));
    defparam add_33905_13.INIT0 = 16'hf555;
    defparam add_33905_13.INIT1 = 16'hf555;
    defparam add_33905_13.INJECT1_0 = "NO";
    defparam add_33905_13.INJECT1_1 = "NO";
    CCU2D add_33905_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48790), .COUT(n48791));
    defparam add_33905_11.INIT0 = 16'hf555;
    defparam add_33905_11.INIT1 = 16'hf555;
    defparam add_33905_11.INJECT1_0 = "NO";
    defparam add_33905_11.INJECT1_1 = "NO";
    CCU2D add_33905_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48789), .COUT(n48790));
    defparam add_33905_9.INIT0 = 16'hf555;
    defparam add_33905_9.INIT1 = 16'hf555;
    defparam add_33905_9.INJECT1_0 = "NO";
    defparam add_33905_9.INJECT1_1 = "NO";
    CCU2D add_33905_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48788), .COUT(n48789));
    defparam add_33905_7.INIT0 = 16'hf555;
    defparam add_33905_7.INIT1 = 16'hf555;
    defparam add_33905_7.INJECT1_0 = "NO";
    defparam add_33905_7.INJECT1_1 = "NO";
    CCU2D add_33905_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48787), .COUT(n48788));
    defparam add_33905_5.INIT0 = 16'hf555;
    defparam add_33905_5.INIT1 = 16'hf555;
    defparam add_33905_5.INJECT1_0 = "NO";
    defparam add_33905_5.INJECT1_1 = "NO";
    CCU2D add_33905_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48786), .COUT(n48787));
    defparam add_33905_3.INIT0 = 16'hf555;
    defparam add_33905_3.INIT1 = 16'hf555;
    defparam add_33905_3.INJECT1_0 = "NO";
    defparam add_33905_3.INJECT1_1 = "NO";
    CCU2D add_33905_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48786));
    defparam add_33905_1.INIT0 = 16'hF000;
    defparam add_33905_1.INIT1 = 16'ha666;
    defparam add_33905_1.INJECT1_0 = "NO";
    defparam add_33905_1.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47699), .COUT(n47700), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47698), .COUT(n47699), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47697), .COUT(n47698), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47696), .COUT(n47697), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47695), .COUT(n47696), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47694), .COUT(n47695), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47693), .COUT(n47694), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47693), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47691), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47690), .COUT(n47691), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_3114_33 (.A0(bit_counter[31]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48322), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_33.INIT0 = 16'h5999;
    defparam add_3114_33.INIT1 = 16'h0000;
    defparam add_3114_33.INJECT1_0 = "NO";
    defparam add_3114_33.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47689), .COUT(n47690), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47688), .COUT(n47689), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_3114_31 (.A0(bit_counter[29]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48321), .COUT(n48322), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_31.INIT0 = 16'h5999;
    defparam add_3114_31.INIT1 = 16'h5999;
    defparam add_3114_31.INJECT1_0 = "NO";
    defparam add_3114_31.INJECT1_1 = "NO";
    CCU2D add_3114_29 (.A0(bit_counter[27]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48320), .COUT(n48321), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_29.INIT0 = 16'h5999;
    defparam add_3114_29.INIT1 = 16'h5999;
    defparam add_3114_29.INJECT1_0 = "NO";
    defparam add_3114_29.INJECT1_1 = "NO";
    CCU2D add_3114_27 (.A0(bit_counter[25]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48319), .COUT(n48320), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_27.INIT0 = 16'h5999;
    defparam add_3114_27.INIT1 = 16'h5999;
    defparam add_3114_27.INJECT1_0 = "NO";
    defparam add_3114_27.INJECT1_1 = "NO";
    CCU2D add_3114_25 (.A0(bit_counter[23]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48318), .COUT(n48319), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_25.INIT0 = 16'h5999;
    defparam add_3114_25.INIT1 = 16'h5999;
    defparam add_3114_25.INJECT1_0 = "NO";
    defparam add_3114_25.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47688), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3114_23 (.A0(bit_counter[21]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48317), .COUT(n48318), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_23.INIT0 = 16'h5999;
    defparam add_3114_23.INIT1 = 16'h5999;
    defparam add_3114_23.INJECT1_0 = "NO";
    defparam add_3114_23.INJECT1_1 = "NO";
    CCU2D add_3114_21 (.A0(bit_counter[19]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48316), .COUT(n48317), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_21.INIT0 = 16'h5999;
    defparam add_3114_21.INIT1 = 16'h5999;
    defparam add_3114_21.INJECT1_0 = "NO";
    defparam add_3114_21.INJECT1_1 = "NO";
    CCU2D add_3114_19 (.A0(bit_counter[17]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48315), .COUT(n48316), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_19.INIT0 = 16'h5999;
    defparam add_3114_19.INIT1 = 16'h5999;
    defparam add_3114_19.INJECT1_0 = "NO";
    defparam add_3114_19.INJECT1_1 = "NO";
    CCU2D add_3114_17 (.A0(bit_counter[15]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48314), .COUT(n48315), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_17.INIT0 = 16'h5999;
    defparam add_3114_17.INIT1 = 16'h5999;
    defparam add_3114_17.INJECT1_0 = "NO";
    defparam add_3114_17.INJECT1_1 = "NO";
    CCU2D add_3114_15 (.A0(bit_counter[13]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48313), .COUT(n48314), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_15.INIT0 = 16'h5999;
    defparam add_3114_15.INIT1 = 16'h5999;
    defparam add_3114_15.INJECT1_0 = "NO";
    defparam add_3114_15.INJECT1_1 = "NO";
    CCU2D add_3114_13 (.A0(bit_counter[11]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48312), .COUT(n48313), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_13.INIT0 = 16'h5999;
    defparam add_3114_13.INIT1 = 16'h5999;
    defparam add_3114_13.INJECT1_0 = "NO";
    defparam add_3114_13.INJECT1_1 = "NO";
    CCU2D add_3114_11 (.A0(bit_counter[9]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48311), .COUT(n48312), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_11.INIT0 = 16'h5999;
    defparam add_3114_11.INIT1 = 16'h5999;
    defparam add_3114_11.INJECT1_0 = "NO";
    defparam add_3114_11.INJECT1_1 = "NO";
    CCU2D add_3114_9 (.A0(bit_counter[7]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48310), .COUT(n48311), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_9.INIT0 = 16'h5999;
    defparam add_3114_9.INIT1 = 16'h5999;
    defparam add_3114_9.INJECT1_0 = "NO";
    defparam add_3114_9.INJECT1_1 = "NO";
    CCU2D add_3114_7 (.A0(bit_counter[5]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48309), .COUT(n48310), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_7.INIT0 = 16'h5999;
    defparam add_3114_7.INIT1 = 16'h5999;
    defparam add_3114_7.INJECT1_0 = "NO";
    defparam add_3114_7.INJECT1_1 = "NO";
    CCU2D add_3114_5 (.A0(bit_counter[3]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48308), .COUT(n48309), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_5.INIT0 = 16'h5999;
    defparam add_3114_5.INIT1 = 16'h5999;
    defparam add_3114_5.INJECT1_0 = "NO";
    defparam add_3114_5.INJECT1_1 = "NO";
    CCU2D add_3114_3 (.A0(bit_counter[1]), .B0(n13276), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13276), .C1(GND_net), 
          .D1(GND_net), .CIN(n48307), .COUT(n48308), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_3.INIT0 = 16'h5999;
    defparam add_3114_3.INIT1 = 16'h5999;
    defparam add_3114_3.INJECT1_0 = "NO";
    defparam add_3114_3.INJECT1_1 = "NO";
    CCU2D add_3114_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13276), .C1(GND_net), .D1(GND_net), 
          .COUT(n48307), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3114_1.INIT0 = 16'hF000;
    defparam add_3114_1.INIT1 = 16'h5999;
    defparam add_3114_1.INJECT1_0 = "NO";
    defparam add_3114_1.INJECT1_1 = "NO";
    PFUMX i38935 (.BLUT(n54940), .ALUT(n54941), .C0(state[1]), .Z(n54942));
    PFUMX i38925 (.BLUT(n54925), .ALUT(n54926), .C0(state[0]), .Z(n54927));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U39 
//

module \WS2812(48000000,"111111111")_U39  (\port_status[0] , sclk_c, ws2813_out_c_0, 
            GND_net, \Q[0] , \RdAddress[0] );
    output \port_status[0] ;
    input sclk_c;
    output ws2813_out_c_0;
    input GND_net;
    input [23:0]\Q[0] ;
    output [8:0]\RdAddress[0] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire sclk_c_enable_11, n54834, sclk_c_enable_12, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_16;
    wire [2:0]state_2__N_104;
    
    wire n47534;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    wire [31:0]n447;
    
    wire n47533, n47532, n47531, n47530, n47529, n47528, n47527, 
        n47526, n47525, n12891, n47524, n47523, n47522, n47521, 
        n47520, n47519, n11271, n54862, n54863, n54864, n47517;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]n118;
    
    wire n47516, n47515, n47514, n54920, n54919, sclk_c_enable_1240, 
        n52935, n53242;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire serial_N_437, n53240, n53241, n54674, n54732, n54731, sclk_c_enable_1241;
    wire [31:0]n6610;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1239, n34738, sclk_c_enable_1238;
    wire [8:0]cur_pixel_8__N_107;
    wire [31:0]bit_counter_31__N_172;
    
    wire n52921, n52922, n52929, n1, n1_adj_904, n52923, n52924, 
        n52930, n52925, n52926, n52931, n15, n14, n42576, n52927, 
        n52928, n52932, n12856, n54617, n103, n34661, n54835;
    wire [31:0]n6434;
    
    wire n76, n34657, n54921, n68, n69;
    wire [6:0]n14998;
    wire [31:0]bit_counter_31__N_204;
    
    wire n39914, n54662, n54608, n52715, n6609, n53239, n53238, 
        n53237, n53236, n52933, n52934, n4, n48402, n48401, n48400, 
        n48399, n48398, n48397, n48396, n48395, n48394, n48393, 
        n48392, n48391, n48390, n48389, n48388, n48387, n48673, 
        n48672, n48671, n48670, n48669, n48668, n48667, n48666, 
        n48665, n48664, n48663, n48662, n48661, n48660, n48659, 
        n48658, n48641, n48640, n48639, n48638, n48637, n48636, 
        n48635, n48634, n48633, n48632, n48631, n48630, n48629, 
        n48628, n48627, n48626;
    
    FD1P3AX status_77 (.D(n54834), .SP(sclk_c_enable_11), .CK(sclk_c), 
            .Q(\port_status[0] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_12), .CK(sclk_c), 
            .Q(ws2813_out_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_16), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_16), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_16), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47534), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47533), .COUT(n47534), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47532), .COUT(n47533), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47531), .COUT(n47532), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47530), .COUT(n47531), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47529), .COUT(n47530), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47528), .COUT(n47529), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47527), .COUT(n47528), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47526), .COUT(n47527), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47525), .COUT(n47526), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    LUT4 i38445_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n12891), .Z(sclk_c_enable_16)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38445_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47524), .COUT(n47525), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47523), .COUT(n47524), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47522), .COUT(n47523), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47521), .COUT(n47522), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47520), .COUT(n47521), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47519), .COUT(n47520), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47519), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n12891), .Z(n11271)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    PFUMX i38883 (.BLUT(n54862), .ALUT(n54863), .C0(state[1]), .Z(n54864));
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47517), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47516), .COUT(n47517), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47515), .COUT(n47516), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47514), .COUT(n47515), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47514), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 mux_2012_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n12891), .Z(n54920)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2012_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2012_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n12891), .Z(n54919)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2012_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 i38404_2_lut_rep_787 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1240)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38404_2_lut_rep_787.init = 16'h9999;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n52935), .B(n53242), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    L6MUX21 i38036 (.D0(n53240), .D1(n53241), .SD(bit_counter[2]), .Z(n53242));
    LUT4 mux_3049_i1_4_lut (.A(n54674), .B(n54732), .C(n11271), .D(n54731), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3049_i1_4_lut.init = 16'h3f3a;
    FD1P3AX delay_counter_i0_i1 (.D(n6610[1]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3IX pixel_i23 (.D(\Q[0] [23]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[0] [22]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[0] [21]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[0] [20]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[0] [19]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[0] [18]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[0] [17]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[0] [16]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[0] [15]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[0] [14]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[0] [13]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[0] [12]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[0] [11]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[0] [10]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[0] [9]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[0] [8]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[0] [7]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[0] [6]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[0] [5]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[0] [4]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[0] [3]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[0] [2]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[0] [1]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n6610[3]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n6610[7]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n6610[8]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n6610[9]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n6610[12]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    PFUMX i37723 (.BLUT(n52921), .ALUT(n52922), .C0(bit_counter[1]), .Z(n52929));
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1240), .CD(n34738), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_904), .SP(sclk_c_enable_1240), .CD(n34738), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    PFUMX i37724 (.BLUT(n52923), .ALUT(n52924), .C0(bit_counter[1]), .Z(n52930));
    PFUMX i37725 (.BLUT(n52925), .ALUT(n52926), .C0(bit_counter[1]), .Z(n52931));
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[7]), .C(n14), .D(cur_pixel[4]), 
         .Z(n42576)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    PFUMX i37726 (.BLUT(n52927), .ALUT(n52928), .C0(bit_counter[1]), .Z(n52932));
    LUT4 i1_2_lut_rep_671 (.A(n42576), .B(n12856), .Z(n54674)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_671.init = 16'h8888;
    LUT4 i1_2_lut_rep_614_3_lut (.A(n42576), .B(n12856), .C(state[1]), 
         .Z(n54617)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_614_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42576), .B(n12856), .C(n54731), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n54617), .B(n54835), .C(n447[7]), .D(n54731), 
         .Z(n6434[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_333 (.A(n54617), .B(n54835), .C(n447[8]), 
         .D(n54731), .Z(n6434[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_333.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_334 (.A(n54617), .B(n54835), .C(n447[9]), 
         .D(n54731), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_334.init = 16'hf888;
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    LUT4 i6_4_lut (.A(cur_pixel[2]), .B(cur_pixel[8]), .C(cur_pixel[6]), 
         .D(cur_pixel[5]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[3]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1241), 
            .CD(n34661), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1241), .CD(n34661), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1241), .CD(n34661), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54921), .SP(sclk_c_enable_1241), .CD(n34657), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54864), .SP(sclk_c_enable_1241), .CD(n34657), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_728_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54731)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_728_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_335 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_335.init = 16'he0f0;
    LUT4 i1_3_lut_rep_708_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1239)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_708_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n14998[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_729_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54732)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_729_3_lut.init = 16'hf8f8;
    LUT4 i22589_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n34738)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22589_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n12891), 
         .Z(sclk_c_enable_12)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i27727_1_lut_rep_831 (.A(state[2]), .Z(n54834)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27727_1_lut_rep_831.init = 16'h5555;
    LUT4 i1_2_lut_3_lut_3_lut (.A(state[2]), .B(bit_counter_31__N_204[15]), 
         .C(state[0]), .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n12856), 
         .D(state[0]), .Z(n39914)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i38479_3_lut_rep_611_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), 
         .D(n12891), .Z(sclk_c_enable_1241)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38479_3_lut_rep_611_4_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_3_lut_3_lut_adj_336 (.A(state[2]), .B(bit_counter_31__N_204[14]), 
         .C(state[0]), .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_336.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_337 (.A(state[2]), .B(bit_counter_31__N_204[13]), 
         .C(state[0]), .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_337.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_338 (.A(state[2]), .B(bit_counter_31__N_204[9]), 
         .C(state[0]), .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_338.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_339 (.A(state[2]), .B(bit_counter_31__N_204[10]), 
         .C(state[0]), .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_339.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_340 (.A(state[2]), .B(bit_counter_31__N_204[21]), 
         .C(state[0]), .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_340.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_341 (.A(state[2]), .B(bit_counter_31__N_204[12]), 
         .C(state[0]), .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_341.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_342 (.A(state[2]), .B(bit_counter_31__N_204[16]), 
         .C(state[0]), .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_342.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_343 (.A(state[2]), .B(bit_counter_31__N_204[11]), 
         .C(state[0]), .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_343.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_344 (.A(state[2]), .B(bit_counter_31__N_204[17]), 
         .C(state[0]), .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_344.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_345 (.A(state[2]), .B(bit_counter_31__N_204[18]), 
         .C(state[0]), .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_345.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_346 (.A(state[2]), .B(bit_counter_31__N_204[31]), 
         .C(state[0]), .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_346.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_347 (.A(state[2]), .B(bit_counter_31__N_204[30]), 
         .C(state[0]), .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_347.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_348 (.A(state[2]), .B(bit_counter_31__N_204[19]), 
         .C(state[0]), .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_348.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_349 (.A(state[2]), .B(bit_counter_31__N_204[29]), 
         .C(state[0]), .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_349.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_350 (.A(state[2]), .B(bit_counter_31__N_204[28]), 
         .C(state[0]), .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_350.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_351 (.A(state[2]), .B(bit_counter_31__N_204[27]), 
         .C(state[0]), .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_351.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_352 (.A(state[2]), .B(bit_counter_31__N_204[26]), 
         .C(state[0]), .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_352.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_353 (.A(state[2]), .B(bit_counter_31__N_204[0]), 
         .C(state[0]), .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_353.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_354 (.A(state[2]), .B(bit_counter_31__N_204[25]), 
         .C(state[0]), .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_354.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_355 (.A(state[2]), .B(bit_counter_31__N_204[24]), 
         .C(state[0]), .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_355.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_356 (.A(state[2]), .B(bit_counter_31__N_204[1]), 
         .C(state[0]), .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_356.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_357 (.A(state[2]), .B(bit_counter_31__N_204[23]), 
         .C(state[0]), .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_357.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_358 (.A(state[2]), .B(bit_counter_31__N_204[20]), 
         .C(state[0]), .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_358.init = 16'h4040;
    LUT4 i1_2_lut_rep_659_2_lut (.A(state[2]), .B(n12891), .Z(n54662)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_659_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_3_lut_adj_359 (.A(state[2]), .B(bit_counter_31__N_204[22]), 
         .C(state[0]), .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_359.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_360 (.A(state[2]), .B(bit_counter_31__N_204[2]), 
         .C(state[0]), .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_360.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_361 (.A(state[2]), .B(bit_counter_31__N_204[5]), 
         .C(state[0]), .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_361.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_362 (.A(state[2]), .B(bit_counter_31__N_204[6]), 
         .C(state[0]), .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_362.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_363 (.A(state[2]), .B(bit_counter_31__N_204[7]), 
         .C(state[0]), .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_363.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_3_lut_adj_364 (.A(state[2]), .B(bit_counter_31__N_204[8]), 
         .C(state[0]), .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_3_lut_adj_364.init = 16'h4040;
    LUT4 i1_2_lut_rep_605_3_lut_3_lut (.A(state[2]), .B(state[1]), .C(n12891), 
         .Z(n54608)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_605_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_365 (.A(state[2]), .B(n42576), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_365.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_366 (.A(state[2]), .B(n42576), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_366.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_367 (.A(state[2]), .B(n42576), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_367.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_368 (.A(state[2]), .B(n42576), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_368.init = 16'h1010;
    LUT4 i28818_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28818_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_2_lut_rep_832 (.A(state[2]), .B(state[0]), .Z(n54835)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_832.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_369 (.A(state[2]), .B(n42576), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_369.init = 16'h1010;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[0]), .C(n12856), 
         .D(state[1]), .Z(sclk_c_enable_1238)) /* synthesis lut_function=(A (D)+!A !(((D)+!C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'haa40;
    LUT4 i1_2_lut_3_lut_adj_370 (.A(state[2]), .B(n42576), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_370.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_371 (.A(state[2]), .B(n42576), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_371.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_372 (.A(state[2]), .B(n42576), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_372.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_373 (.A(state[2]), .B(n42576), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_373.init = 16'h1010;
    FD1P3IX pixel_i0 (.D(\Q[0] [0]), .SP(sclk_c_enable_1239), .CD(n34738), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1238), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1239), 
            .CD(n34738), .CK(sclk_c), .Q(\RdAddress[0] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1240), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i0 (.D(n6610[0]), .SP(sclk_c_enable_1241), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=135, LSE_RLINE=135 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54835), .B(state[1]), .C(n54674), .D(n54662), 
         .Z(n52715)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 mux_3049_i2_4_lut_4_lut (.A(n54732), .B(n54731), .C(n11271), 
         .D(n12856), .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_3049_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 mux_2022_i2_4_lut (.A(n68), .B(n14998[0]), .C(n6609), .D(n52715), 
         .Z(n6610[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i2_4_lut.init = 16'hcfca;
    LUT4 i2034_3_lut (.A(state[2]), .B(state[1]), .C(n12891), .Z(n6609)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2034_3_lut.init = 16'ha8a8;
    LUT4 i38033_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38033_3_lut.init = 16'hcaca;
    LUT4 i38032_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38032_3_lut.init = 16'hcaca;
    LUT4 i38031_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38031_3_lut.init = 16'hcaca;
    LUT4 i38030_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53236)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38030_3_lut.init = 16'hcaca;
    LUT4 mux_2022_i1_4_lut (.A(n69), .B(n14998[0]), .C(n6609), .D(n52715), 
         .Z(n6610[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i1_4_lut.init = 16'hcfca;
    L6MUX21 i37729 (.D0(n52933), .D1(n52934), .SD(bit_counter[3]), .Z(n52935));
    PFUMX i38034 (.BLUT(n53236), .ALUT(n53237), .C0(bit_counter[1]), .Z(n53240));
    PFUMX i38035 (.BLUT(n53238), .ALUT(n53239), .C0(bit_counter[1]), .Z(n53241));
    L6MUX21 i37727 (.D0(n52929), .D1(n52930), .SD(bit_counter[2]), .Z(n52933));
    L6MUX21 i37728 (.D0(n52931), .D1(n52932), .SD(bit_counter[2]), .Z(n52934));
    LUT4 mux_2022_i4_4_lut (.A(n39914), .B(n54732), .C(n6609), .D(n4), 
         .Z(n6610[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42576), .B(n54608), .C(n447[3]), .D(n54731), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2022_i8_4_lut (.A(n6434[7]), .B(n54732), .C(n6609), .D(n54608), 
         .Z(n6610[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i8_4_lut.init = 16'h303a;
    LUT4 mux_2022_i9_4_lut (.A(n6434[8]), .B(n54732), .C(n6609), .D(n54608), 
         .Z(n6610[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i9_4_lut.init = 16'h303a;
    LUT4 mux_2022_i10_4_lut (.A(n76), .B(n54732), .C(n6609), .D(n54608), 
         .Z(n6610[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i10_4_lut.init = 16'h303a;
    LUT4 mux_2022_i13_4_lut (.A(n54608), .B(n54732), .C(n6609), .D(n103), 
         .Z(n6610[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2022_i13_4_lut.init = 16'h3530;
    LUT4 i37722_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n52928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37722_3_lut.init = 16'hcaca;
    LUT4 i37721_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n52927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37721_3_lut.init = 16'hcaca;
    LUT4 i37720_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n52926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37720_3_lut.init = 16'hcaca;
    LUT4 i37719_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n52925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37719_3_lut.init = 16'hcaca;
    LUT4 i37718_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37718_3_lut.init = 16'hcaca;
    LUT4 i37717_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37717_3_lut.init = 16'hcaca;
    LUT4 i37716_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37716_3_lut.init = 16'hcaca;
    LUT4 i37715_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37715_3_lut.init = 16'hcaca;
    LUT4 i28762_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28762_2_lut.init = 16'hbbbb;
    LUT4 i28763_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_904)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28763_2_lut.init = 16'hbbbb;
    LUT4 i22445_2_lut_4_lut (.A(n54662), .B(state[0]), .C(state[1]), .D(n6609), 
         .Z(n34657)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i22445_2_lut_4_lut.init = 16'hfd00;
    CCU2D add_3102_33 (.A0(bit_counter[31]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48402), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_33.INIT0 = 16'h5999;
    defparam add_3102_33.INIT1 = 16'h0000;
    defparam add_3102_33.INJECT1_0 = "NO";
    defparam add_3102_33.INJECT1_1 = "NO";
    CCU2D add_3102_31 (.A0(bit_counter[29]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48401), .COUT(n48402), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_31.INIT0 = 16'h5999;
    defparam add_3102_31.INIT1 = 16'h5999;
    defparam add_3102_31.INJECT1_0 = "NO";
    defparam add_3102_31.INJECT1_1 = "NO";
    CCU2D add_3102_29 (.A0(bit_counter[27]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48400), .COUT(n48401), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_29.INIT0 = 16'h5999;
    defparam add_3102_29.INIT1 = 16'h5999;
    defparam add_3102_29.INJECT1_0 = "NO";
    defparam add_3102_29.INJECT1_1 = "NO";
    CCU2D add_3102_27 (.A0(bit_counter[25]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48399), .COUT(n48400), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_27.INIT0 = 16'h5999;
    defparam add_3102_27.INIT1 = 16'h5999;
    defparam add_3102_27.INJECT1_0 = "NO";
    defparam add_3102_27.INJECT1_1 = "NO";
    LUT4 i22469_4_lut (.A(sclk_c_enable_1241), .B(n54731), .C(n6609), 
         .D(n54608), .Z(n34661)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22469_4_lut.init = 16'haaa2;
    CCU2D add_3102_25 (.A0(bit_counter[23]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48398), .COUT(n48399), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_25.INIT0 = 16'h5999;
    defparam add_3102_25.INIT1 = 16'h5999;
    defparam add_3102_25.INJECT1_0 = "NO";
    defparam add_3102_25.INJECT1_1 = "NO";
    CCU2D add_3102_23 (.A0(bit_counter[21]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48397), .COUT(n48398), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_23.INIT0 = 16'h5999;
    defparam add_3102_23.INIT1 = 16'h5999;
    defparam add_3102_23.INJECT1_0 = "NO";
    defparam add_3102_23.INJECT1_1 = "NO";
    CCU2D add_3102_21 (.A0(bit_counter[19]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48396), .COUT(n48397), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_21.INIT0 = 16'h5999;
    defparam add_3102_21.INIT1 = 16'h5999;
    defparam add_3102_21.INJECT1_0 = "NO";
    defparam add_3102_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54674), .C(n12891), .D(n54835), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    CCU2D add_3102_19 (.A0(bit_counter[17]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48395), .COUT(n48396), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_19.INIT0 = 16'h5999;
    defparam add_3102_19.INIT1 = 16'h5999;
    defparam add_3102_19.INJECT1_0 = "NO";
    defparam add_3102_19.INJECT1_1 = "NO";
    CCU2D add_3102_17 (.A0(bit_counter[15]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48394), .COUT(n48395), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_17.INIT0 = 16'h5999;
    defparam add_3102_17.INIT1 = 16'h5999;
    defparam add_3102_17.INJECT1_0 = "NO";
    defparam add_3102_17.INJECT1_1 = "NO";
    CCU2D add_3102_15 (.A0(bit_counter[13]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48393), .COUT(n48394), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_15.INIT0 = 16'h5999;
    defparam add_3102_15.INIT1 = 16'h5999;
    defparam add_3102_15.INJECT1_0 = "NO";
    defparam add_3102_15.INJECT1_1 = "NO";
    CCU2D add_3102_13 (.A0(bit_counter[11]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48392), .COUT(n48393), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_13.INIT0 = 16'h5999;
    defparam add_3102_13.INIT1 = 16'h5999;
    defparam add_3102_13.INJECT1_0 = "NO";
    defparam add_3102_13.INJECT1_1 = "NO";
    CCU2D add_3102_11 (.A0(bit_counter[9]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48391), .COUT(n48392), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_11.INIT0 = 16'h5999;
    defparam add_3102_11.INIT1 = 16'h5999;
    defparam add_3102_11.INJECT1_0 = "NO";
    defparam add_3102_11.INJECT1_1 = "NO";
    CCU2D add_3102_9 (.A0(bit_counter[7]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48390), .COUT(n48391), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_9.INIT0 = 16'h5999;
    defparam add_3102_9.INIT1 = 16'h5999;
    defparam add_3102_9.INJECT1_0 = "NO";
    defparam add_3102_9.INJECT1_1 = "NO";
    CCU2D add_3102_7 (.A0(bit_counter[5]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48389), .COUT(n48390), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_7.INIT0 = 16'h5999;
    defparam add_3102_7.INIT1 = 16'h5999;
    defparam add_3102_7.INJECT1_0 = "NO";
    defparam add_3102_7.INJECT1_1 = "NO";
    CCU2D add_3102_5 (.A0(bit_counter[3]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48388), .COUT(n48389), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_5.INIT0 = 16'h5999;
    defparam add_3102_5.INIT1 = 16'h5999;
    defparam add_3102_5.INJECT1_0 = "NO";
    defparam add_3102_5.INJECT1_1 = "NO";
    CCU2D add_3102_3 (.A0(bit_counter[1]), .B0(n12856), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n12856), .C1(GND_net), 
          .D1(GND_net), .CIN(n48387), .COUT(n48388), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_3.INIT0 = 16'h5999;
    defparam add_3102_3.INIT1 = 16'h5999;
    defparam add_3102_3.INJECT1_0 = "NO";
    defparam add_3102_3.INJECT1_1 = "NO";
    CCU2D add_3102_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n12856), .C1(GND_net), .D1(GND_net), 
          .COUT(n48387), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3102_1.INIT0 = 16'hF000;
    defparam add_3102_1.INIT1 = 16'h5999;
    defparam add_3102_1.INJECT1_0 = "NO";
    defparam add_3102_1.INJECT1_1 = "NO";
    LUT4 mux_2012_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n12891), .Z(n54863)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2012_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2012_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n12856), .Z(n54862)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2012_i3_4_lut_else_4_lut.init = 16'hd0f2;
    CCU2D add_33942_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48673), 
          .S0(n12891));
    defparam add_33942_cout.INIT0 = 16'h0000;
    defparam add_33942_cout.INIT1 = 16'h0000;
    defparam add_33942_cout.INJECT1_0 = "NO";
    defparam add_33942_cout.INJECT1_1 = "NO";
    CCU2D add_33942_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48672), .COUT(n48673));
    defparam add_33942_31.INIT0 = 16'hf555;
    defparam add_33942_31.INIT1 = 16'h5555;
    defparam add_33942_31.INJECT1_0 = "NO";
    defparam add_33942_31.INJECT1_1 = "NO";
    CCU2D add_33942_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48671), .COUT(n48672));
    defparam add_33942_29.INIT0 = 16'hf555;
    defparam add_33942_29.INIT1 = 16'hf555;
    defparam add_33942_29.INJECT1_0 = "NO";
    defparam add_33942_29.INJECT1_1 = "NO";
    CCU2D add_33942_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48670), .COUT(n48671));
    defparam add_33942_27.INIT0 = 16'hf555;
    defparam add_33942_27.INIT1 = 16'hf555;
    defparam add_33942_27.INJECT1_0 = "NO";
    defparam add_33942_27.INJECT1_1 = "NO";
    CCU2D add_33942_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48669), .COUT(n48670));
    defparam add_33942_25.INIT0 = 16'hf555;
    defparam add_33942_25.INIT1 = 16'hf555;
    defparam add_33942_25.INJECT1_0 = "NO";
    defparam add_33942_25.INJECT1_1 = "NO";
    CCU2D add_33942_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48668), .COUT(n48669));
    defparam add_33942_23.INIT0 = 16'hf555;
    defparam add_33942_23.INIT1 = 16'hf555;
    defparam add_33942_23.INJECT1_0 = "NO";
    defparam add_33942_23.INJECT1_1 = "NO";
    CCU2D add_33942_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48667), .COUT(n48668));
    defparam add_33942_21.INIT0 = 16'hf555;
    defparam add_33942_21.INIT1 = 16'hf555;
    defparam add_33942_21.INJECT1_0 = "NO";
    defparam add_33942_21.INJECT1_1 = "NO";
    CCU2D add_33942_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48666), .COUT(n48667));
    defparam add_33942_19.INIT0 = 16'hf555;
    defparam add_33942_19.INIT1 = 16'hf555;
    defparam add_33942_19.INJECT1_0 = "NO";
    defparam add_33942_19.INJECT1_1 = "NO";
    CCU2D add_33942_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48665), .COUT(n48666));
    defparam add_33942_17.INIT0 = 16'hf555;
    defparam add_33942_17.INIT1 = 16'hf555;
    defparam add_33942_17.INJECT1_0 = "NO";
    defparam add_33942_17.INJECT1_1 = "NO";
    CCU2D add_33942_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48664), .COUT(n48665));
    defparam add_33942_15.INIT0 = 16'hf555;
    defparam add_33942_15.INIT1 = 16'hf555;
    defparam add_33942_15.INJECT1_0 = "NO";
    defparam add_33942_15.INJECT1_1 = "NO";
    CCU2D add_33942_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48663), .COUT(n48664));
    defparam add_33942_13.INIT0 = 16'hf555;
    defparam add_33942_13.INIT1 = 16'hf555;
    defparam add_33942_13.INJECT1_0 = "NO";
    defparam add_33942_13.INJECT1_1 = "NO";
    CCU2D add_33942_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48662), .COUT(n48663));
    defparam add_33942_11.INIT0 = 16'hf555;
    defparam add_33942_11.INIT1 = 16'hf555;
    defparam add_33942_11.INJECT1_0 = "NO";
    defparam add_33942_11.INJECT1_1 = "NO";
    CCU2D add_33942_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48661), .COUT(n48662));
    defparam add_33942_9.INIT0 = 16'hf555;
    defparam add_33942_9.INIT1 = 16'hf555;
    defparam add_33942_9.INJECT1_0 = "NO";
    defparam add_33942_9.INJECT1_1 = "NO";
    CCU2D add_33942_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48660), .COUT(n48661));
    defparam add_33942_7.INIT0 = 16'hf555;
    defparam add_33942_7.INIT1 = 16'hf555;
    defparam add_33942_7.INJECT1_0 = "NO";
    defparam add_33942_7.INJECT1_1 = "NO";
    CCU2D add_33942_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48659), .COUT(n48660));
    defparam add_33942_5.INIT0 = 16'hf555;
    defparam add_33942_5.INIT1 = 16'hf555;
    defparam add_33942_5.INJECT1_0 = "NO";
    defparam add_33942_5.INJECT1_1 = "NO";
    CCU2D add_33942_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48658), .COUT(n48659));
    defparam add_33942_3.INIT0 = 16'hf555;
    defparam add_33942_3.INIT1 = 16'hf555;
    defparam add_33942_3.INJECT1_0 = "NO";
    defparam add_33942_3.INJECT1_1 = "NO";
    CCU2D add_33942_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48658));
    defparam add_33942_1.INIT0 = 16'hF000;
    defparam add_33942_1.INIT1 = 16'ha666;
    defparam add_33942_1.INJECT1_0 = "NO";
    defparam add_33942_1.INJECT1_1 = "NO";
    CCU2D add_33943_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48641), 
          .S0(n12856));
    defparam add_33943_cout.INIT0 = 16'h0000;
    defparam add_33943_cout.INIT1 = 16'h0000;
    defparam add_33943_cout.INJECT1_0 = "NO";
    defparam add_33943_cout.INJECT1_1 = "NO";
    CCU2D add_33943_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48640), .COUT(n48641));
    defparam add_33943_31.INIT0 = 16'hf555;
    defparam add_33943_31.INIT1 = 16'h5555;
    defparam add_33943_31.INJECT1_0 = "NO";
    defparam add_33943_31.INJECT1_1 = "NO";
    CCU2D add_33943_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48639), .COUT(n48640));
    defparam add_33943_29.INIT0 = 16'hf555;
    defparam add_33943_29.INIT1 = 16'hf555;
    defparam add_33943_29.INJECT1_0 = "NO";
    defparam add_33943_29.INJECT1_1 = "NO";
    CCU2D add_33943_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48638), .COUT(n48639));
    defparam add_33943_27.INIT0 = 16'hf555;
    defparam add_33943_27.INIT1 = 16'hf555;
    defparam add_33943_27.INJECT1_0 = "NO";
    defparam add_33943_27.INJECT1_1 = "NO";
    CCU2D add_33943_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48637), .COUT(n48638));
    defparam add_33943_25.INIT0 = 16'hf555;
    defparam add_33943_25.INIT1 = 16'hf555;
    defparam add_33943_25.INJECT1_0 = "NO";
    defparam add_33943_25.INJECT1_1 = "NO";
    CCU2D add_33943_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48636), .COUT(n48637));
    defparam add_33943_23.INIT0 = 16'hf555;
    defparam add_33943_23.INIT1 = 16'hf555;
    defparam add_33943_23.INJECT1_0 = "NO";
    defparam add_33943_23.INJECT1_1 = "NO";
    CCU2D add_33943_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48635), .COUT(n48636));
    defparam add_33943_21.INIT0 = 16'hf555;
    defparam add_33943_21.INIT1 = 16'hf555;
    defparam add_33943_21.INJECT1_0 = "NO";
    defparam add_33943_21.INJECT1_1 = "NO";
    CCU2D add_33943_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48634), .COUT(n48635));
    defparam add_33943_19.INIT0 = 16'hf555;
    defparam add_33943_19.INIT1 = 16'hf555;
    defparam add_33943_19.INJECT1_0 = "NO";
    defparam add_33943_19.INJECT1_1 = "NO";
    CCU2D add_33943_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48633), .COUT(n48634));
    defparam add_33943_17.INIT0 = 16'hf555;
    defparam add_33943_17.INIT1 = 16'hf555;
    defparam add_33943_17.INJECT1_0 = "NO";
    defparam add_33943_17.INJECT1_1 = "NO";
    CCU2D add_33943_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48632), .COUT(n48633));
    defparam add_33943_15.INIT0 = 16'hf555;
    defparam add_33943_15.INIT1 = 16'hf555;
    defparam add_33943_15.INJECT1_0 = "NO";
    defparam add_33943_15.INJECT1_1 = "NO";
    CCU2D add_33943_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48631), .COUT(n48632));
    defparam add_33943_13.INIT0 = 16'hf555;
    defparam add_33943_13.INIT1 = 16'hf555;
    defparam add_33943_13.INJECT1_0 = "NO";
    defparam add_33943_13.INJECT1_1 = "NO";
    CCU2D add_33943_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48630), .COUT(n48631));
    defparam add_33943_11.INIT0 = 16'hf555;
    defparam add_33943_11.INIT1 = 16'hf555;
    defparam add_33943_11.INJECT1_0 = "NO";
    defparam add_33943_11.INJECT1_1 = "NO";
    CCU2D add_33943_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48629), .COUT(n48630));
    defparam add_33943_9.INIT0 = 16'hf555;
    defparam add_33943_9.INIT1 = 16'hf555;
    defparam add_33943_9.INJECT1_0 = "NO";
    defparam add_33943_9.INJECT1_1 = "NO";
    CCU2D add_33943_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48628), .COUT(n48629));
    defparam add_33943_7.INIT0 = 16'hf555;
    defparam add_33943_7.INIT1 = 16'hf555;
    defparam add_33943_7.INJECT1_0 = "NO";
    defparam add_33943_7.INJECT1_1 = "NO";
    CCU2D add_33943_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48627), .COUT(n48628));
    defparam add_33943_5.INIT0 = 16'hf555;
    defparam add_33943_5.INIT1 = 16'hf555;
    defparam add_33943_5.INJECT1_0 = "NO";
    defparam add_33943_5.INJECT1_1 = "NO";
    CCU2D add_33943_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48626), .COUT(n48627));
    defparam add_33943_3.INIT0 = 16'hf555;
    defparam add_33943_3.INIT1 = 16'hf555;
    defparam add_33943_3.INJECT1_0 = "NO";
    defparam add_33943_3.INJECT1_1 = "NO";
    CCU2D add_33943_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48626));
    defparam add_33943_1.INIT0 = 16'hF000;
    defparam add_33943_1.INIT1 = 16'ha666;
    defparam add_33943_1.INJECT1_0 = "NO";
    defparam add_33943_1.INJECT1_1 = "NO";
    PFUMX i38921 (.BLUT(n54919), .ALUT(n54920), .C0(state[0]), .Z(n54921));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U28 
//

module \WS2812(48000000,"111111111")_U28  (sclk_c, GND_net, \port_status[1] , 
            ws2813_out_c_1, \Q[1] , \RdAddress[1] );
    input sclk_c;
    input GND_net;
    output \port_status[1] ;
    output ws2813_out_c_1;
    input [23:0]\Q[1] ;
    output [8:0]\RdAddress[1] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_967;
    wire [31:0]n7945;
    
    wire n47558;
    wire [31:0]n447;
    
    wire n47559, n47557, n47556, n47554;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]n118;
    
    wire sclk_c_enable_19, n54816, sclk_c_enable_20, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_24;
    wire [2:0]state_2__N_104;
    
    wire n47553, n47552, n47551, n12961, n12926, sclk_c_enable_1228, 
        n11004, n53247, n53248;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53249, sclk_c_enable_1236, n39746, n54659, n54603, n54689, 
        n15;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1235, n34833;
    wire [8:0]cur_pixel_8__N_107;
    wire [31:0]bit_counter_31__N_172;
    
    wire n1, n1_adj_902, n52944, n52945, n52948, n52946, n52947, 
        n52949, n54810, n34686, serial_N_437, n54843;
    wire [31:0]n7769;
    
    wire n54875, n7944;
    wire [31:0]n7871;
    
    wire n54876, n54874, n52942, n52943, n54720, n58;
    wire [31:0]bit_counter_31__N_204;
    
    wire n52936, n52937;
    wire [6:0]n15040;
    
    wire n52938, n52939, n39779, n39797, n39774, n54557, n52950, 
        n52941, n52940, n53246, n53245, n53244, n53243, n47571, 
        n47570, n47569, n47568, n47567, n47566, n47565, n52636, 
        n47564, n47563, n47562, n47561, n47560, n48386, n48385, 
        n48384, n48383, n48382, n48381, n48380, n48379, n48378, 
        n48377, n48376, n48375, n48374, n48373, n48372, n48371, 
        n15_adj_903, n14, n48737, n48736, n48735, n48734, n48733, 
        n48732, n48731, n48730, n48729, n48728, n48727, n48726, 
        n48725, n48724, n48723, n48722, n48705, n48704, n48703, 
        n48702, n48701, n48700, n48699, n48698, n48697, n48696, 
        n48695, n48694, n48693, n48692, n48691, n48690;
    
    FD1P3AX delay_counter_i0_i0 (.D(n7945[0]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47558), .COUT(n47559), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47557), .COUT(n47558), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47556), .COUT(n47557), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47556), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47554), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    FD1P3AX status_77 (.D(n54816), .SP(sclk_c_enable_19), .CK(sclk_c), 
            .Q(\port_status[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_20), .CK(sclk_c), 
            .Q(ws2813_out_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_24), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_24), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_24), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47553), .COUT(n47554), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47552), .COUT(n47553), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47551), .COUT(n47552), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47551), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i38633_3_lut_rep_567_4_lut (.A(state[2]), .B(n12961), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_967)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38633_3_lut_rep_567_4_lut.init = 16'hfffb;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n12926), 
         .D(state[0]), .Z(sclk_c_enable_1228)) /* synthesis lut_function=(A (B)+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h9888;
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n12961), .Z(n11004)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 i2_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n12961), 
         .D(state[0]), .Z(sclk_c_enable_24)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_4_lut.init = 16'hf9f8;
    L6MUX21 i38043 (.D0(n53247), .D1(n53248), .SD(bit_counter[2]), .Z(n53249));
    LUT4 i38412_2_lut_rep_792 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1236)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38412_2_lut_rep_792.init = 16'h9999;
    LUT4 i1_2_lut_rep_656 (.A(n12926), .B(n39746), .Z(n54659)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_656.init = 16'h8888;
    LUT4 i1_2_lut_rep_600_3_lut (.A(n12926), .B(n39746), .C(state[1]), 
         .Z(n54603)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_600_3_lut.init = 16'h0808;
    LUT4 i29482_3_lut_4_lut (.A(n12926), .B(n39746), .C(n54689), .D(n447[12]), 
         .Z(n15)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i29482_3_lut_4_lut.init = 16'hf808;
    FD1P3IX pixel_i23 (.D(\Q[1] [23]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[1] [22]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[1] [21]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[1] [20]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[1] [19]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[1] [18]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[1] [17]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[1] [16]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[1] [15]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[1] [14]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[1] [13]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[1] [12]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[1] [11]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[1] [10]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[1] [9]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[1] [8]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[1] [7]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[1] [6]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[1] [5]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[1] [4]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[1] [3]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[1] [2]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[1] [1]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1236), .CD(n34833), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_902), .SP(sclk_c_enable_1236), .CD(n34833), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i1 (.D(n7945[1]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n7945[3]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n7945[7]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n7945[8]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n7945[9]), .SP(sclk_c_enable_967), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n7945[12]), .SP(sclk_c_enable_967), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    L6MUX21 i37742 (.D0(n52944), .D1(n52945), .SD(bit_counter[2]), .Z(n52948));
    L6MUX21 i37743 (.D0(n52946), .D1(n52947), .SD(bit_counter[2]), .Z(n52949));
    LUT4 i1_2_lut_rep_807 (.A(state[1]), .B(state[2]), .Z(n54810)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_807.init = 16'heeee;
    LUT4 i1_2_lut_rep_686_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54689)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_686_3_lut.init = 16'hefef;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    LUT4 i27637_1_lut_rep_813 (.A(state[2]), .Z(n54816)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i27637_1_lut_rep_813.init = 16'h5555;
    LUT4 i28823_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28823_3_lut_3_lut.init = 16'h5151;
    LUT4 i2_3_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[7]), .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2_3_lut_3_lut.init = 16'h1010;
    LUT4 i1_3_lut_4_lut (.A(n54603), .B(n54843), .C(n447[7]), .D(n54689), 
         .Z(n7769[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_301 (.A(n54603), .B(n54843), .C(n447[8]), 
         .D(n54689), .Z(n7769[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_301.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_302 (.A(n54603), .B(n54843), .C(n447[9]), 
         .D(n54689), .Z(n7769[9])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_302.init = 16'hf888;
    LUT4 mux_2297_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n12961), .Z(n54875)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2297_i3_4_lut_then_4_lut.init = 16'hd1f0;
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_967), 
            .CD(n34686), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_967), .CD(n34686), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_967), .CD(n34686), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n7871[4]), .SP(sclk_c_enable_967), .CD(n7944), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54876), .SP(sclk_c_enable_967), .CD(n7944), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 mux_2297_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n12926), .Z(n54874)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2297_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i30059_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[8]), .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i30059_2_lut_3_lut.init = 16'h1010;
    LUT4 i29428_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[6]), .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29428_2_lut_3_lut.init = 16'h1010;
    LUT4 i29427_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[5]), .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29427_2_lut_3_lut.init = 16'h1010;
    LUT4 i29426_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[4]), .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29426_2_lut_3_lut.init = 16'h1010;
    LUT4 i29425_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[3]), .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29425_2_lut_3_lut.init = 16'h1010;
    LUT4 i29424_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[2]), .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29424_2_lut_3_lut.init = 16'h1010;
    LUT4 i29423_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[1]), .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29423_2_lut_3_lut.init = 16'h1010;
    LUT4 i28821_2_lut_3_lut (.A(state[2]), .B(n39746), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i28821_2_lut_3_lut.init = 16'h1010;
    FD1P3IX pixel_i0 (.D(\Q[1] [0]), .SP(sclk_c_enable_1235), .CD(n34833), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1228), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1235), 
            .CD(n34833), .CK(sclk_c), .Q(\RdAddress[1] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1236), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=146, LSE_RLINE=146 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    PFUMX i37741 (.BLUT(n52942), .ALUT(n52943), .C0(bit_counter[1]), .Z(n52947));
    LUT4 mux_2992_i2_4_lut_4_lut (.A(n54720), .B(n54689), .C(n11004), 
         .D(n12926), .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2992_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_840 (.A(state[0]), .B(state[2]), .Z(n54843)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_840.init = 16'h2222;
    LUT4 i2_2_lut_3_lut_4_lut (.A(state[0]), .B(state[2]), .C(n12926), 
         .D(state[1]), .Z(n58)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    PFUMX i37738 (.BLUT(n52936), .ALUT(n52937), .C0(bit_counter[1]), .Z(n52944));
    LUT4 i1_2_lut_3_lut_adj_303 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_303.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_304 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_304.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_305 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_305.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_306 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_306.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_307 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_307.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_308 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_308.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_309 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_309.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_310 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_310.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_311 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_311.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_312 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_312.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_313 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_313.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_314 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_314.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_315 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_315.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_316 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_316.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_317 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_317.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_318 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_318.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_319 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_319.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_320 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_320.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_321 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_321.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_322 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_322.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_323 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_323.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_324 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_324.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_325 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_325.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_326 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_326.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_327 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_327.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_328 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_328.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_329 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_329.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_330 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_330.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_331 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_331.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n12961), 
         .Z(sclk_c_enable_20)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i22684_2_lut_4_lut_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n34833)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22684_2_lut_4_lut_2_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_717_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54720)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_717_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_adj_332 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15040[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_332.init = 16'h7070;
    LUT4 i1_3_lut_rep_710_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1235)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i1_3_lut_rep_710_4_lut_3_lut.init = 16'h8989;
    PFUMX i37739 (.BLUT(n52938), .ALUT(n52939), .C0(bit_counter[1]), .Z(n52945));
    LUT4 i29490_3_lut_4_lut (.A(state[0]), .B(n54810), .C(n447[0]), .D(n39746), 
         .Z(n39779)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29490_3_lut_4_lut.init = 16'hd0f2;
    LUT4 i29494_3_lut_4_lut (.A(state[0]), .B(n54810), .C(n447[1]), .D(n39746), 
         .Z(n39797)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29494_3_lut_4_lut.init = 16'hd0f2;
    LUT4 i29486_3_lut_4_lut (.A(state[0]), .B(n54810), .C(n447[3]), .D(n39746), 
         .Z(n39774)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29486_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_2297_i5_4_lut_4_lut (.A(state[0]), .B(n54810), .C(n447[4]), 
         .D(n54557), .Z(n7871[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2297_i5_4_lut_4_lut.init = 16'haad0;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n52950), .B(n53249), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i37735_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n52941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37735_3_lut.init = 16'hcaca;
    LUT4 i37734_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n52940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37734_3_lut.init = 16'hcaca;
    LUT4 i38040_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38040_3_lut.init = 16'hcaca;
    LUT4 i38039_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38039_3_lut.init = 16'hcaca;
    LUT4 i38038_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38038_3_lut.init = 16'hcaca;
    LUT4 i38037_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38037_3_lut.init = 16'hcaca;
    LUT4 mux_2992_i1_4_lut (.A(n54659), .B(n54720), .C(n11004), .D(n54689), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2992_i1_4_lut.init = 16'h3f3a;
    LUT4 i37733_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n52939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37733_3_lut.init = 16'hcaca;
    LUT4 i37732_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n52938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37732_3_lut.init = 16'hcaca;
    LUT4 i37731_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n52937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37731_3_lut.init = 16'hcaca;
    LUT4 i37730_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n52936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37730_3_lut.init = 16'hcaca;
    PFUMX i38041 (.BLUT(n53243), .ALUT(n53244), .C0(bit_counter[1]), .Z(n53247));
    PFUMX i38042 (.BLUT(n53245), .ALUT(n53246), .C0(bit_counter[1]), .Z(n53248));
    PFUMX i37740 (.BLUT(n52940), .ALUT(n52941), .C0(bit_counter[1]), .Z(n52946));
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47571), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    L6MUX21 i37744 (.D0(n52948), .D1(n52949), .SD(bit_counter[3]), .Z(n52950));
    LUT4 i37737_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n52943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37737_3_lut.init = 16'hcaca;
    LUT4 i37736_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n52942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37736_3_lut.init = 16'hcaca;
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47570), .COUT(n47571), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47569), .COUT(n47570), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47568), .COUT(n47569), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47567), .COUT(n47568), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    LUT4 i28758_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28758_2_lut.init = 16'hbbbb;
    LUT4 i28761_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_902)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28761_2_lut.init = 16'hbbbb;
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47566), .COUT(n47567), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47565), .COUT(n47566), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    LUT4 mux_2307_i2_4_lut (.A(n39797), .B(n15040[0]), .C(n7944), .D(n52636), 
         .Z(n7945[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2307_i4_4_lut (.A(n39774), .B(n54720), .C(n7944), .D(n52636), 
         .Z(n7945[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i4_4_lut.init = 16'h3f3a;
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47564), .COUT(n47565), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    LUT4 mux_2307_i8_4_lut (.A(n7769[7]), .B(n54720), .C(n7944), .D(n54557), 
         .Z(n7945[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i8_4_lut.init = 16'h303a;
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47563), .COUT(n47564), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    LUT4 mux_2307_i9_4_lut (.A(n7769[8]), .B(n54720), .C(n7944), .D(n54557), 
         .Z(n7945[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i9_4_lut.init = 16'h303a;
    PFUMX i38891 (.BLUT(n54874), .ALUT(n54875), .C0(state[1]), .Z(n54876));
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47562), .COUT(n47563), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    LUT4 mux_2307_i10_4_lut (.A(n7769[9]), .B(n54720), .C(n7944), .D(n54557), 
         .Z(n7945[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i10_4_lut.init = 16'h303a;
    LUT4 mux_2307_i13_4_lut (.A(n54557), .B(n54720), .C(n7944), .D(n15), 
         .Z(n7945[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i13_4_lut.init = 16'h3530;
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47561), .COUT(n47562), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47560), .COUT(n47561), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47559), .COUT(n47560), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54659), .C(n12961), .D(n54843), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    LUT4 i22494_4_lut (.A(sclk_c_enable_967), .B(n54689), .C(n7944), .D(n54557), 
         .Z(n34686)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i22494_4_lut.init = 16'haaa2;
    CCU2D add_3104_33 (.A0(bit_counter[31]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48386), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_33.INIT0 = 16'h5999;
    defparam add_3104_33.INIT1 = 16'h0000;
    defparam add_3104_33.INJECT1_0 = "NO";
    defparam add_3104_33.INJECT1_1 = "NO";
    CCU2D add_3104_31 (.A0(bit_counter[29]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48385), .COUT(n48386), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_31.INIT0 = 16'h5999;
    defparam add_3104_31.INIT1 = 16'h5999;
    defparam add_3104_31.INJECT1_0 = "NO";
    defparam add_3104_31.INJECT1_1 = "NO";
    CCU2D add_3104_29 (.A0(bit_counter[27]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48384), .COUT(n48385), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_29.INIT0 = 16'h5999;
    defparam add_3104_29.INIT1 = 16'h5999;
    defparam add_3104_29.INJECT1_0 = "NO";
    defparam add_3104_29.INJECT1_1 = "NO";
    CCU2D add_3104_27 (.A0(bit_counter[25]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48383), .COUT(n48384), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_27.INIT0 = 16'h5999;
    defparam add_3104_27.INIT1 = 16'h5999;
    defparam add_3104_27.INJECT1_0 = "NO";
    defparam add_3104_27.INJECT1_1 = "NO";
    CCU2D add_3104_25 (.A0(bit_counter[23]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48382), .COUT(n48383), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_25.INIT0 = 16'h5999;
    defparam add_3104_25.INIT1 = 16'h5999;
    defparam add_3104_25.INJECT1_0 = "NO";
    defparam add_3104_25.INJECT1_1 = "NO";
    CCU2D add_3104_23 (.A0(bit_counter[21]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48381), .COUT(n48382), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_23.INIT0 = 16'h5999;
    defparam add_3104_23.INIT1 = 16'h5999;
    defparam add_3104_23.INJECT1_0 = "NO";
    defparam add_3104_23.INJECT1_1 = "NO";
    CCU2D add_3104_21 (.A0(bit_counter[19]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48380), .COUT(n48381), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_21.INIT0 = 16'h5999;
    defparam add_3104_21.INIT1 = 16'h5999;
    defparam add_3104_21.INJECT1_0 = "NO";
    defparam add_3104_21.INJECT1_1 = "NO";
    CCU2D add_3104_19 (.A0(bit_counter[17]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48379), .COUT(n48380), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_19.INIT0 = 16'h5999;
    defparam add_3104_19.INIT1 = 16'h5999;
    defparam add_3104_19.INJECT1_0 = "NO";
    defparam add_3104_19.INJECT1_1 = "NO";
    CCU2D add_3104_17 (.A0(bit_counter[15]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48378), .COUT(n48379), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_17.INIT0 = 16'h5999;
    defparam add_3104_17.INIT1 = 16'h5999;
    defparam add_3104_17.INJECT1_0 = "NO";
    defparam add_3104_17.INJECT1_1 = "NO";
    CCU2D add_3104_15 (.A0(bit_counter[13]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48377), .COUT(n48378), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_15.INIT0 = 16'h5999;
    defparam add_3104_15.INIT1 = 16'h5999;
    defparam add_3104_15.INJECT1_0 = "NO";
    defparam add_3104_15.INJECT1_1 = "NO";
    CCU2D add_3104_13 (.A0(bit_counter[11]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48376), .COUT(n48377), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_13.INIT0 = 16'h5999;
    defparam add_3104_13.INIT1 = 16'h5999;
    defparam add_3104_13.INJECT1_0 = "NO";
    defparam add_3104_13.INJECT1_1 = "NO";
    LUT4 mux_2307_i1_4_lut (.A(n39779), .B(n15040[0]), .C(n7944), .D(n52636), 
         .Z(n7945[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2307_i1_4_lut.init = 16'hcfca;
    CCU2D add_3104_11 (.A0(bit_counter[9]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48375), .COUT(n48376), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_11.INIT0 = 16'h5999;
    defparam add_3104_11.INIT1 = 16'h5999;
    defparam add_3104_11.INJECT1_0 = "NO";
    defparam add_3104_11.INJECT1_1 = "NO";
    CCU2D add_3104_9 (.A0(bit_counter[7]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48374), .COUT(n48375), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_9.INIT0 = 16'h5999;
    defparam add_3104_9.INIT1 = 16'h5999;
    defparam add_3104_9.INJECT1_0 = "NO";
    defparam add_3104_9.INJECT1_1 = "NO";
    CCU2D add_3104_7 (.A0(bit_counter[5]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48373), .COUT(n48374), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_7.INIT0 = 16'h5999;
    defparam add_3104_7.INIT1 = 16'h5999;
    defparam add_3104_7.INJECT1_0 = "NO";
    defparam add_3104_7.INJECT1_1 = "NO";
    CCU2D add_3104_5 (.A0(bit_counter[3]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48372), .COUT(n48373), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_5.INIT0 = 16'h5999;
    defparam add_3104_5.INIT1 = 16'h5999;
    defparam add_3104_5.INJECT1_0 = "NO";
    defparam add_3104_5.INJECT1_1 = "NO";
    CCU2D add_3104_3 (.A0(bit_counter[1]), .B0(n12926), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n12926), .C1(GND_net), 
          .D1(GND_net), .CIN(n48371), .COUT(n48372), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_3.INIT0 = 16'h5999;
    defparam add_3104_3.INIT1 = 16'h5999;
    defparam add_3104_3.INJECT1_0 = "NO";
    defparam add_3104_3.INJECT1_1 = "NO";
    CCU2D add_3104_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n12926), .C1(GND_net), .D1(GND_net), 
          .COUT(n48371), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3104_1.INIT0 = 16'hF000;
    defparam add_3104_1.INIT1 = 16'h5999;
    defparam add_3104_1.INJECT1_0 = "NO";
    defparam add_3104_1.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n15_adj_903), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[2]), 
         .Z(n39746)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[8]), .B(cur_pixel[7]), .C(cur_pixel[1]), 
         .D(cur_pixel[6]), .Z(n15_adj_903)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[5]), .B(cur_pixel[0]), .C(cur_pixel[3]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i5_3_lut.init = 16'h8080;
    CCU2D add_33939_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48737), 
          .S0(n12961));
    defparam add_33939_cout.INIT0 = 16'h0000;
    defparam add_33939_cout.INIT1 = 16'h0000;
    defparam add_33939_cout.INJECT1_0 = "NO";
    defparam add_33939_cout.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[2]), .B(n12961), .C(n58), .D(state[1]), 
         .Z(n52636)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf4f0;
    CCU2D add_33939_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48736), .COUT(n48737));
    defparam add_33939_31.INIT0 = 16'hf555;
    defparam add_33939_31.INIT1 = 16'h5555;
    defparam add_33939_31.INJECT1_0 = "NO";
    defparam add_33939_31.INJECT1_1 = "NO";
    CCU2D add_33939_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48735), .COUT(n48736));
    defparam add_33939_29.INIT0 = 16'hf555;
    defparam add_33939_29.INIT1 = 16'hf555;
    defparam add_33939_29.INJECT1_0 = "NO";
    defparam add_33939_29.INJECT1_1 = "NO";
    CCU2D add_33939_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48734), .COUT(n48735));
    defparam add_33939_27.INIT0 = 16'hf555;
    defparam add_33939_27.INIT1 = 16'hf555;
    defparam add_33939_27.INJECT1_0 = "NO";
    defparam add_33939_27.INJECT1_1 = "NO";
    CCU2D add_33939_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48733), .COUT(n48734));
    defparam add_33939_25.INIT0 = 16'hf555;
    defparam add_33939_25.INIT1 = 16'hf555;
    defparam add_33939_25.INJECT1_0 = "NO";
    defparam add_33939_25.INJECT1_1 = "NO";
    CCU2D add_33939_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48732), .COUT(n48733));
    defparam add_33939_23.INIT0 = 16'hf555;
    defparam add_33939_23.INIT1 = 16'hf555;
    defparam add_33939_23.INJECT1_0 = "NO";
    defparam add_33939_23.INJECT1_1 = "NO";
    CCU2D add_33939_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48731), .COUT(n48732));
    defparam add_33939_21.INIT0 = 16'hf555;
    defparam add_33939_21.INIT1 = 16'hf555;
    defparam add_33939_21.INJECT1_0 = "NO";
    defparam add_33939_21.INJECT1_1 = "NO";
    CCU2D add_33939_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48730), .COUT(n48731));
    defparam add_33939_19.INIT0 = 16'hf555;
    defparam add_33939_19.INIT1 = 16'hf555;
    defparam add_33939_19.INJECT1_0 = "NO";
    defparam add_33939_19.INJECT1_1 = "NO";
    CCU2D add_33939_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48729), .COUT(n48730));
    defparam add_33939_17.INIT0 = 16'hf555;
    defparam add_33939_17.INIT1 = 16'hf555;
    defparam add_33939_17.INJECT1_0 = "NO";
    defparam add_33939_17.INJECT1_1 = "NO";
    CCU2D add_33939_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48728), .COUT(n48729));
    defparam add_33939_15.INIT0 = 16'hf555;
    defparam add_33939_15.INIT1 = 16'hf555;
    defparam add_33939_15.INJECT1_0 = "NO";
    defparam add_33939_15.INJECT1_1 = "NO";
    CCU2D add_33939_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48727), .COUT(n48728));
    defparam add_33939_13.INIT0 = 16'hf555;
    defparam add_33939_13.INIT1 = 16'hf555;
    defparam add_33939_13.INJECT1_0 = "NO";
    defparam add_33939_13.INJECT1_1 = "NO";
    CCU2D add_33939_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48726), .COUT(n48727));
    defparam add_33939_11.INIT0 = 16'hf555;
    defparam add_33939_11.INIT1 = 16'hf555;
    defparam add_33939_11.INJECT1_0 = "NO";
    defparam add_33939_11.INJECT1_1 = "NO";
    CCU2D add_33939_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48725), .COUT(n48726));
    defparam add_33939_9.INIT0 = 16'hf555;
    defparam add_33939_9.INIT1 = 16'hf555;
    defparam add_33939_9.INJECT1_0 = "NO";
    defparam add_33939_9.INJECT1_1 = "NO";
    CCU2D add_33939_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48724), .COUT(n48725));
    defparam add_33939_7.INIT0 = 16'hf555;
    defparam add_33939_7.INIT1 = 16'hf555;
    defparam add_33939_7.INJECT1_0 = "NO";
    defparam add_33939_7.INJECT1_1 = "NO";
    CCU2D add_33939_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48723), .COUT(n48724));
    defparam add_33939_5.INIT0 = 16'hf555;
    defparam add_33939_5.INIT1 = 16'hf555;
    defparam add_33939_5.INJECT1_0 = "NO";
    defparam add_33939_5.INJECT1_1 = "NO";
    CCU2D add_33939_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48722), .COUT(n48723));
    defparam add_33939_3.INIT0 = 16'hf555;
    defparam add_33939_3.INIT1 = 16'hf555;
    defparam add_33939_3.INJECT1_0 = "NO";
    defparam add_33939_3.INJECT1_1 = "NO";
    CCU2D add_33939_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48722));
    defparam add_33939_1.INIT0 = 16'hF000;
    defparam add_33939_1.INIT1 = 16'ha666;
    defparam add_33939_1.INJECT1_0 = "NO";
    defparam add_33939_1.INJECT1_1 = "NO";
    CCU2D add_33941_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48705), 
          .S0(n12926));
    defparam add_33941_cout.INIT0 = 16'h0000;
    defparam add_33941_cout.INIT1 = 16'h0000;
    defparam add_33941_cout.INJECT1_0 = "NO";
    defparam add_33941_cout.INJECT1_1 = "NO";
    CCU2D add_33941_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48704), .COUT(n48705));
    defparam add_33941_31.INIT0 = 16'hf555;
    defparam add_33941_31.INIT1 = 16'h5555;
    defparam add_33941_31.INJECT1_0 = "NO";
    defparam add_33941_31.INJECT1_1 = "NO";
    CCU2D add_33941_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48703), .COUT(n48704));
    defparam add_33941_29.INIT0 = 16'hf555;
    defparam add_33941_29.INIT1 = 16'hf555;
    defparam add_33941_29.INJECT1_0 = "NO";
    defparam add_33941_29.INJECT1_1 = "NO";
    CCU2D add_33941_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48702), .COUT(n48703));
    defparam add_33941_27.INIT0 = 16'hf555;
    defparam add_33941_27.INIT1 = 16'hf555;
    defparam add_33941_27.INJECT1_0 = "NO";
    defparam add_33941_27.INJECT1_1 = "NO";
    CCU2D add_33941_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48701), .COUT(n48702));
    defparam add_33941_25.INIT0 = 16'hf555;
    defparam add_33941_25.INIT1 = 16'hf555;
    defparam add_33941_25.INJECT1_0 = "NO";
    defparam add_33941_25.INJECT1_1 = "NO";
    CCU2D add_33941_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48700), .COUT(n48701));
    defparam add_33941_23.INIT0 = 16'hf555;
    defparam add_33941_23.INIT1 = 16'hf555;
    defparam add_33941_23.INJECT1_0 = "NO";
    defparam add_33941_23.INJECT1_1 = "NO";
    CCU2D add_33941_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48699), .COUT(n48700));
    defparam add_33941_21.INIT0 = 16'hf555;
    defparam add_33941_21.INIT1 = 16'hf555;
    defparam add_33941_21.INJECT1_0 = "NO";
    defparam add_33941_21.INJECT1_1 = "NO";
    CCU2D add_33941_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48698), .COUT(n48699));
    defparam add_33941_19.INIT0 = 16'hf555;
    defparam add_33941_19.INIT1 = 16'hf555;
    defparam add_33941_19.INJECT1_0 = "NO";
    defparam add_33941_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_554_3_lut (.A(state[2]), .B(n12961), .C(state[1]), 
         .Z(n54557)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_554_3_lut.init = 16'h4040;
    CCU2D add_33941_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48697), .COUT(n48698));
    defparam add_33941_17.INIT0 = 16'hf555;
    defparam add_33941_17.INIT1 = 16'hf555;
    defparam add_33941_17.INJECT1_0 = "NO";
    defparam add_33941_17.INJECT1_1 = "NO";
    CCU2D add_33941_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48696), .COUT(n48697));
    defparam add_33941_15.INIT0 = 16'hf555;
    defparam add_33941_15.INIT1 = 16'hf555;
    defparam add_33941_15.INJECT1_0 = "NO";
    defparam add_33941_15.INJECT1_1 = "NO";
    CCU2D add_33941_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48695), .COUT(n48696));
    defparam add_33941_13.INIT0 = 16'hf555;
    defparam add_33941_13.INIT1 = 16'hf555;
    defparam add_33941_13.INJECT1_0 = "NO";
    defparam add_33941_13.INJECT1_1 = "NO";
    CCU2D add_33941_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48694), .COUT(n48695));
    defparam add_33941_11.INIT0 = 16'hf555;
    defparam add_33941_11.INIT1 = 16'hf555;
    defparam add_33941_11.INJECT1_0 = "NO";
    defparam add_33941_11.INJECT1_1 = "NO";
    CCU2D add_33941_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48693), .COUT(n48694));
    defparam add_33941_9.INIT0 = 16'hf555;
    defparam add_33941_9.INIT1 = 16'hf555;
    defparam add_33941_9.INJECT1_0 = "NO";
    defparam add_33941_9.INJECT1_1 = "NO";
    CCU2D add_33941_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48692), .COUT(n48693));
    defparam add_33941_7.INIT0 = 16'hf555;
    defparam add_33941_7.INIT1 = 16'hf555;
    defparam add_33941_7.INJECT1_0 = "NO";
    defparam add_33941_7.INJECT1_1 = "NO";
    CCU2D add_33941_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48691), .COUT(n48692));
    defparam add_33941_5.INIT0 = 16'hf555;
    defparam add_33941_5.INIT1 = 16'hf555;
    defparam add_33941_5.INJECT1_0 = "NO";
    defparam add_33941_5.INJECT1_1 = "NO";
    CCU2D add_33941_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48690), .COUT(n48691));
    defparam add_33941_3.INIT0 = 16'hf555;
    defparam add_33941_3.INIT1 = 16'hf555;
    defparam add_33941_3.INJECT1_0 = "NO";
    defparam add_33941_3.INJECT1_1 = "NO";
    CCU2D add_33941_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48690));
    defparam add_33941_1.INIT0 = 16'hF000;
    defparam add_33941_1.INIT1 = 16'ha666;
    defparam add_33941_1.INJECT1_0 = "NO";
    defparam add_33941_1.INJECT1_1 = "NO";
    LUT4 i2319_3_lut (.A(state[2]), .B(state[1]), .C(n12961), .Z(n7944)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2319_3_lut.init = 16'ha8a8;
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U32 
//

module \WS2812(48000000,"111111111")_U32  (sclk_c, \port_status[16] , ws2813_out_c_16, 
            \Q[16] , \RdAddress[16] , GND_net);
    input sclk_c;
    output \port_status[16] ;
    output ws2813_out_c_16;
    input [23:0]\Q[16] ;
    output [8:0]\RdAddress[16] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    wire [31:0]bit_counter_31__N_204;
    wire [31:0]bit_counter_31__N_172;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1840;
    wire [31:0]n10126;
    
    wire sclk_c_enable_146, n54763, sclk_c_enable_147, serial_N_433, 
        sclk_c_enable_151;
    wire [2:0]state_2__N_104;
    
    wire n54865, n54866, n54867, n42684, n13976, n54638, n14011, 
        n54569, n53169, n53170;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53173, n54639, n54580, n53171, n53172, n53174;
    wire [31:0]n447;
    
    wire n71;
    wire [6:0]n15105;
    
    wire n10125, n52667, n37883, n41613, n4, n54704;
    wire [31:0]n9950;
    
    wire n80, n53352, n53353, n53354, n54774;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1658, n36258;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire sclk_c_enable_1625;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1689, n54868;
    wire [8:0]n118;
    
    wire n48545, n48544, n48543, n48542, n48541, n48540, n53161, 
        n53162, n53163, n53164, n53165, n53166, n53167, n53168, 
        n53351, n53350, n53349, n53348, n48539, n36076, n54775;
    wire [31:0]n10052;
    wire [2:0]n7204;
    
    wire n48538, n48537, n48536, n48535, n48534, n48533, n48532, 
        n48531, n48530, n74, n53175, n48513, n48512, n48511, n48510, 
        n48509, n48508, n48507, n48506, n48505, n48504, n48503, 
        n48502, n48501, n48500, n48499, n48498, n36229, n1, n1_adj_901, 
        n36080, n54869, n47951, n47950, n47949, n47948, n47947, 
        n47946, n47945, n47944, n47943, n47942, n47941, n47940, 
        n47939, n47938, n47937, n47936, n15, n14, serial_N_437, 
        n54631, n7211, n48062, n48061, n48060, n48059, n48058, 
        n48057, n48056, n48055, n48054, n48053, n48052, n48051, 
        n48050, n48049, n48048, n48047, n48045, n48044, n48043, 
        n48042;
    
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_254 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_254.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_255 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_255.init = 16'h2020;
    FD1P3AX delay_counter_i0_i0 (.D(n10126[0]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54763), .SP(sclk_c_enable_146), .CK(sclk_c), 
            .Q(\port_status[16] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_147), .CK(sclk_c), 
            .Q(ws2813_out_c_16)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_151), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_151), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_151), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    PFUMX i38885 (.BLUT(n54865), .ALUT(n54866), .C0(state[1]), .Z(n54867));
    LUT4 i1_2_lut_3_lut_adj_256 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_256.init = 16'h2020;
    LUT4 i1_2_lut_rep_635 (.A(n42684), .B(n13976), .Z(n54638)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_635.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n14011), .Z(sclk_c_enable_151)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i1_2_lut_rep_566_3_lut (.A(n42684), .B(n13976), .C(state[1]), 
         .Z(n54569)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_566_3_lut.init = 16'h0808;
    L6MUX21 i37967 (.D0(n53169), .D1(n53170), .SD(bit_counter[2]), .Z(n53173));
    LUT4 i1_2_lut_rep_636 (.A(state[2]), .B(n14011), .Z(n54639)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_636.init = 16'h4444;
    LUT4 i1_2_lut_rep_577_3_lut (.A(state[2]), .B(n14011), .C(state[1]), 
         .Z(n54580)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_577_3_lut.init = 16'h4040;
    LUT4 i38578_3_lut_rep_578_4_lut (.A(state[2]), .B(n14011), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1840)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i38578_3_lut_rep_578_4_lut.init = 16'hfffb;
    L6MUX21 i37968 (.D0(n53171), .D1(n53172), .SD(bit_counter[2]), .Z(n53174));
    LUT4 mux_2780_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14011), .Z(n54866)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2780_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2790_i2_4_lut (.A(n71), .B(n15105[0]), .C(n10125), .D(n52667), 
         .Z(n10126[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2790_i4_4_lut (.A(n37883), .B(n41613), .C(n10125), .D(n4), 
         .Z(n10126[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n42684), .B(n54580), .C(n447[3]), .D(n54704), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 i1_2_lut_3_lut_adj_257 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_257.init = 16'h2020;
    LUT4 mux_2790_i8_4_lut (.A(n9950[7]), .B(n41613), .C(n10125), .D(n54580), 
         .Z(n10126[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i8_4_lut.init = 16'h303a;
    LUT4 i1_2_lut_3_lut_adj_258 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_258.init = 16'h2020;
    LUT4 mux_2790_i9_4_lut (.A(n9950[8]), .B(n41613), .C(n10125), .D(n54580), 
         .Z(n10126[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i9_4_lut.init = 16'h303a;
    LUT4 mux_2780_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13976), .Z(n54865)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2780_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 mux_2790_i10_4_lut (.A(n80), .B(n41613), .C(n10125), .D(n54580), 
         .Z(n10126[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i10_4_lut.init = 16'h303a;
    LUT4 mux_2790_i13_4_lut (.A(n9950[12]), .B(n41613), .C(n10125), .D(n54580), 
         .Z(n10126[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i13_4_lut.init = 16'h303a;
    LUT4 i1_2_lut_3_lut_adj_259 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15105[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_259.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_adj_260 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_260.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_261 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_261.init = 16'h2020;
    L6MUX21 i38148 (.D0(n53352), .D1(n53353), .SD(bit_counter[2]), .Z(n53354));
    LUT4 i29444_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n41613)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i29444_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_771 (.A(state[0]), .B(state[2]), .Z(n54774)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_771.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_262 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_262.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_263 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_263.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13976), 
         .D(state[1]), .Z(n37883)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_adj_264 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_264.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_265 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_265.init = 16'h2020;
    FD1P3IX pixel_i0 (.D(\Q[16] [0]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13976), 
         .D(state[1]), .Z(sclk_c_enable_1625)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_266 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_266.init = 16'h2020;
    LUT4 i38566_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n13976), 
         .Z(n54868)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38566_4_lut_else_3_lut.init = 16'h0404;
    FD1P3AX delay_counter_i0_i1 (.D(n10126[1]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n10126[3]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n10126[7]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n10126[8]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n10126[9]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n10126[12]), .SP(sclk_c_enable_1840), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_267 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_267.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_268 (.A(state[2]), .B(n42684), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_268.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_269 (.A(state[2]), .B(n42684), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_269.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_270 (.A(state[2]), .B(n42684), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_270.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_271 (.A(state[2]), .B(n42684), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_271.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_272 (.A(state[2]), .B(n42684), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_272.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_273 (.A(state[2]), .B(n42684), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_273.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_274 (.A(state[2]), .B(n42684), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_274.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_275 (.A(state[2]), .B(n42684), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_275.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_276 (.A(state[2]), .B(n42684), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_276.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_277 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_277.init = 16'h2020;
    LUT4 i1_3_lut_4_lut (.A(n54569), .B(n54774), .C(n447[8]), .D(n54704), 
         .Z(n9950[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_278 (.A(n54569), .B(n54774), .C(n447[12]), 
         .D(n54704), .Z(n9950[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_278.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_279 (.A(n54569), .B(n54774), .C(n447[9]), 
         .D(n54704), .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_279.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_280 (.A(n54569), .B(n54774), .C(n447[7]), 
         .D(n54704), .Z(n9950[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_280.init = 16'hf888;
    LUT4 i1_2_lut_3_lut_adj_281 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_281.init = 16'h2020;
    CCU2D add_33897_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48545), 
          .S0(n14011));
    defparam add_33897_cout.INIT0 = 16'h0000;
    defparam add_33897_cout.INIT1 = 16'h0000;
    defparam add_33897_cout.INJECT1_0 = "NO";
    defparam add_33897_cout.INJECT1_1 = "NO";
    CCU2D add_33897_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48544), .COUT(n48545));
    defparam add_33897_31.INIT0 = 16'hf555;
    defparam add_33897_31.INIT1 = 16'h5555;
    defparam add_33897_31.INJECT1_0 = "NO";
    defparam add_33897_31.INJECT1_1 = "NO";
    CCU2D add_33897_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48543), .COUT(n48544));
    defparam add_33897_29.INIT0 = 16'hf555;
    defparam add_33897_29.INIT1 = 16'hf555;
    defparam add_33897_29.INJECT1_0 = "NO";
    defparam add_33897_29.INJECT1_1 = "NO";
    CCU2D add_33897_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48542), .COUT(n48543));
    defparam add_33897_27.INIT0 = 16'hf555;
    defparam add_33897_27.INIT1 = 16'hf555;
    defparam add_33897_27.INJECT1_0 = "NO";
    defparam add_33897_27.INJECT1_1 = "NO";
    CCU2D add_33897_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48541), .COUT(n48542));
    defparam add_33897_25.INIT0 = 16'hf555;
    defparam add_33897_25.INIT1 = 16'hf555;
    defparam add_33897_25.INJECT1_0 = "NO";
    defparam add_33897_25.INJECT1_1 = "NO";
    CCU2D add_33897_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48540), .COUT(n48541));
    defparam add_33897_23.INIT0 = 16'hf555;
    defparam add_33897_23.INIT1 = 16'hf555;
    defparam add_33897_23.INJECT1_0 = "NO";
    defparam add_33897_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_282 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_282.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_283 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_283.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_284 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_284.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_285 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_285.init = 16'h2020;
    PFUMX i37963 (.BLUT(n53161), .ALUT(n53162), .C0(bit_counter[1]), .Z(n53169));
    PFUMX i37964 (.BLUT(n53163), .ALUT(n53164), .C0(bit_counter[1]), .Z(n53170));
    LUT4 i1_2_lut_3_lut_adj_286 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_286.init = 16'h2020;
    PFUMX i37965 (.BLUT(n53165), .ALUT(n53166), .C0(bit_counter[1]), .Z(n53171));
    PFUMX i37966 (.BLUT(n53167), .ALUT(n53168), .C0(bit_counter[1]), .Z(n53172));
    LUT4 i38145_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38145_3_lut.init = 16'hcaca;
    LUT4 i38144_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38144_3_lut.init = 16'hcaca;
    LUT4 i38143_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38143_3_lut.init = 16'hcaca;
    LUT4 i38142_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38142_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_287 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_287.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_288 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_288.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_289 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_289.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_290 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_290.init = 16'h2020;
    CCU2D add_33897_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48539), .COUT(n48540));
    defparam add_33897_21.INIT0 = 16'hf555;
    defparam add_33897_21.INIT1 = 16'hf555;
    defparam add_33897_21.INJECT1_0 = "NO";
    defparam add_33897_21.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54774), .B(state[1]), .C(n54638), .D(n54639), 
         .Z(n52667)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 i23864_2_lut_4_lut (.A(n54639), .B(state[0]), .C(state[1]), .D(n10125), 
         .Z(n36076)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23864_2_lut_4_lut.init = 16'hfd00;
    LUT4 mux_2780_i5_4_lut_4_lut (.A(state[0]), .B(n54775), .C(n447[4]), 
         .D(n54580), .Z(n10052[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2780_i5_4_lut_4_lut.init = 16'haad0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_291 (.A(state[0]), .B(n54775), .C(n13976), 
         .D(n42684), .Z(n7204[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_291.init = 16'hfddd;
    LUT4 i1_2_lut_3_lut_adj_292 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_292.init = 16'h2020;
    CCU2D add_33897_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48538), .COUT(n48539));
    defparam add_33897_19.INIT0 = 16'hf555;
    defparam add_33897_19.INIT1 = 16'hf555;
    defparam add_33897_19.INJECT1_0 = "NO";
    defparam add_33897_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_293 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_293.init = 16'h2020;
    CCU2D add_33897_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48537), .COUT(n48538));
    defparam add_33897_17.INIT0 = 16'hf555;
    defparam add_33897_17.INIT1 = 16'hf555;
    defparam add_33897_17.INJECT1_0 = "NO";
    defparam add_33897_17.INJECT1_1 = "NO";
    CCU2D add_33897_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48536), .COUT(n48537));
    defparam add_33897_15.INIT0 = 16'hf555;
    defparam add_33897_15.INIT1 = 16'hf555;
    defparam add_33897_15.INJECT1_0 = "NO";
    defparam add_33897_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_772 (.A(state[1]), .B(state[2]), .Z(n54775)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_772.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_294 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_294.init = 16'h2020;
    CCU2D add_33897_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48535), .COUT(n48536));
    defparam add_33897_13.INIT0 = 16'hf555;
    defparam add_33897_13.INIT1 = 16'hf555;
    defparam add_33897_13.INJECT1_0 = "NO";
    defparam add_33897_13.INJECT1_1 = "NO";
    LUT4 i37962_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37962_3_lut.init = 16'hcaca;
    LUT4 i37961_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37961_3_lut.init = 16'hcaca;
    LUT4 i37960_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37960_3_lut.init = 16'hcaca;
    LUT4 i37959_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37959_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_295 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_295.init = 16'h2020;
    LUT4 i37958_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37958_3_lut.init = 16'hcaca;
    CCU2D add_33897_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48534), .COUT(n48535));
    defparam add_33897_11.INIT0 = 16'hf555;
    defparam add_33897_11.INIT1 = 16'hf555;
    defparam add_33897_11.INJECT1_0 = "NO";
    defparam add_33897_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_296 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_296.init = 16'h2020;
    CCU2D add_33897_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48533), .COUT(n48534));
    defparam add_33897_9.INIT0 = 16'hf555;
    defparam add_33897_9.INIT1 = 16'hf555;
    defparam add_33897_9.INJECT1_0 = "NO";
    defparam add_33897_9.INJECT1_1 = "NO";
    LUT4 i37957_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37957_3_lut.init = 16'hcaca;
    LUT4 i37956_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37956_3_lut.init = 16'hcaca;
    LUT4 i37955_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37955_3_lut.init = 16'hcaca;
    CCU2D add_33897_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48532), .COUT(n48533));
    defparam add_33897_7.INIT0 = 16'hf555;
    defparam add_33897_7.INIT1 = 16'hf555;
    defparam add_33897_7.INJECT1_0 = "NO";
    defparam add_33897_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_701_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54704)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_701_3_lut.init = 16'hefef;
    CCU2D add_33897_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48531), .COUT(n48532));
    defparam add_33897_5.INIT0 = 16'hf555;
    defparam add_33897_5.INIT1 = 16'hf555;
    defparam add_33897_5.INJECT1_0 = "NO";
    defparam add_33897_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n14011), 
         .Z(sclk_c_enable_147)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    CCU2D add_33897_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48530), .COUT(n48531));
    defparam add_33897_3.INIT0 = 16'hf555;
    defparam add_33897_3.INIT1 = 16'hf555;
    defparam add_33897_3.INJECT1_0 = "NO";
    defparam add_33897_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_685_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_1658)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_685_4_lut_3_lut.init = 16'h8989;
    CCU2D add_33897_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48530));
    defparam add_33897_1.INIT0 = 16'hF000;
    defparam add_33897_1.INIT1 = 16'ha666;
    defparam add_33897_1.INJECT1_0 = "NO";
    defparam add_33897_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_297 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_297.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_298 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_298.init = 16'he0f0;
    L6MUX21 i37969 (.D0(n53173), .D1(n53174), .SD(bit_counter[3]), .Z(n53175));
    CCU2D add_33899_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48513), 
          .S0(n13976));
    defparam add_33899_cout.INIT0 = 16'h0000;
    defparam add_33899_cout.INIT1 = 16'h0000;
    defparam add_33899_cout.INJECT1_0 = "NO";
    defparam add_33899_cout.INJECT1_1 = "NO";
    CCU2D add_33899_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48512), .COUT(n48513));
    defparam add_33899_31.INIT0 = 16'hf555;
    defparam add_33899_31.INIT1 = 16'h5555;
    defparam add_33899_31.INJECT1_0 = "NO";
    defparam add_33899_31.INJECT1_1 = "NO";
    CCU2D add_33899_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48511), .COUT(n48512));
    defparam add_33899_29.INIT0 = 16'hf555;
    defparam add_33899_29.INIT1 = 16'hf555;
    defparam add_33899_29.INJECT1_0 = "NO";
    defparam add_33899_29.INJECT1_1 = "NO";
    CCU2D add_33899_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48510), .COUT(n48511));
    defparam add_33899_27.INIT0 = 16'hf555;
    defparam add_33899_27.INIT1 = 16'hf555;
    defparam add_33899_27.INJECT1_0 = "NO";
    defparam add_33899_27.INJECT1_1 = "NO";
    CCU2D add_33899_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48509), .COUT(n48510));
    defparam add_33899_25.INIT0 = 16'hf555;
    defparam add_33899_25.INIT1 = 16'hf555;
    defparam add_33899_25.INJECT1_0 = "NO";
    defparam add_33899_25.INJECT1_1 = "NO";
    CCU2D add_33899_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48508), .COUT(n48509));
    defparam add_33899_23.INIT0 = 16'hf555;
    defparam add_33899_23.INIT1 = 16'hf555;
    defparam add_33899_23.INJECT1_0 = "NO";
    defparam add_33899_23.INJECT1_1 = "NO";
    FD1P3IX pixel_i23 (.D(\Q[16] [23]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[16] [22]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[16] [21]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[16] [20]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[16] [19]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[16] [18]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[16] [17]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[16] [16]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[16] [15]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[16] [14]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[16] [13]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[16] [12]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[16] [11]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[16] [10]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    CCU2D add_33899_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48507), .COUT(n48508));
    defparam add_33899_21.INIT0 = 16'hf555;
    defparam add_33899_21.INIT1 = 16'hf555;
    defparam add_33899_21.INJECT1_0 = "NO";
    defparam add_33899_21.INJECT1_1 = "NO";
    FD1P3IX pixel_i9 (.D(\Q[16] [9]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[16] [8]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[16] [7]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[16] [6]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[16] [5]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[16] [4]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[16] [3]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[16] [2]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[16] [1]), .SP(sclk_c_enable_1658), .CD(n36258), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    PFUMX i38146 (.BLUT(n53348), .ALUT(n53349), .C0(bit_counter[1]), .Z(n53352));
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    PFUMX i38147 (.BLUT(n53350), .ALUT(n53351), .C0(bit_counter[1]), .Z(n53353));
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1625), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    CCU2D add_33899_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48506), .COUT(n48507));
    defparam add_33899_19.INIT0 = 16'hf555;
    defparam add_33899_19.INIT1 = 16'hf555;
    defparam add_33899_19.INJECT1_0 = "NO";
    defparam add_33899_19.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    CCU2D add_33899_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48505), .COUT(n48506));
    defparam add_33899_17.INIT0 = 16'hf555;
    defparam add_33899_17.INIT1 = 16'hf555;
    defparam add_33899_17.INJECT1_0 = "NO";
    defparam add_33899_17.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    CCU2D add_33899_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48504), .COUT(n48505));
    defparam add_33899_15.INIT0 = 16'hf555;
    defparam add_33899_15.INIT1 = 16'hf555;
    defparam add_33899_15.INJECT1_0 = "NO";
    defparam add_33899_15.INJECT1_1 = "NO";
    LUT4 i24109_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n36258)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i24109_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    CCU2D add_33899_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48503), .COUT(n48504));
    defparam add_33899_13.INIT0 = 16'hf555;
    defparam add_33899_13.INIT1 = 16'hf555;
    defparam add_33899_13.INJECT1_0 = "NO";
    defparam add_33899_13.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    CCU2D add_33899_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48502), .COUT(n48503));
    defparam add_33899_11.INIT0 = 16'hf555;
    defparam add_33899_11.INIT1 = 16'hf555;
    defparam add_33899_11.INJECT1_0 = "NO";
    defparam add_33899_11.INJECT1_1 = "NO";
    CCU2D add_33899_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48501), .COUT(n48502));
    defparam add_33899_9.INIT0 = 16'hf555;
    defparam add_33899_9.INIT1 = 16'hf555;
    defparam add_33899_9.INJECT1_0 = "NO";
    defparam add_33899_9.INJECT1_1 = "NO";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1658), 
            .CD(n36258), .CK(sclk_c), .Q(\RdAddress[16] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    CCU2D add_33899_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48500), .COUT(n48501));
    defparam add_33899_7.INIT0 = 16'hf555;
    defparam add_33899_7.INIT1 = 16'hf555;
    defparam add_33899_7.INJECT1_0 = "NO";
    defparam add_33899_7.INJECT1_1 = "NO";
    CCU2D add_33899_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48499), .COUT(n48500));
    defparam add_33899_5.INIT0 = 16'hf555;
    defparam add_33899_5.INIT1 = 16'hf555;
    defparam add_33899_5.INJECT1_0 = "NO";
    defparam add_33899_5.INJECT1_1 = "NO";
    CCU2D add_33899_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48498), .COUT(n48499));
    defparam add_33899_3.INIT0 = 16'hf555;
    defparam add_33899_3.INIT1 = 16'hf555;
    defparam add_33899_3.INJECT1_0 = "NO";
    defparam add_33899_3.INJECT1_1 = "NO";
    CCU2D add_33899_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48498));
    defparam add_33899_1.INIT0 = 16'hF000;
    defparam add_33899_1.INIT1 = 16'ha666;
    defparam add_33899_1.INJECT1_0 = "NO";
    defparam add_33899_1.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1689), .CD(n36229), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_901), .SP(sclk_c_enable_1689), .CD(n36229), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1689), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 i38424_2_lut_rep_746 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1689)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38424_2_lut_rep_746.init = 16'h9999;
    LUT4 i24017_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36229)) /* synthesis lut_function=(A (B)) */ ;
    defparam i24017_2_lut_2_lut.init = 16'h8888;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1840), 
            .CD(n36080), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1840), .CD(n36080), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1840), .CD(n36080), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n10052[4]), .SP(sclk_c_enable_1840), 
            .CD(n36076), .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54867), .SP(sclk_c_enable_1840), .CD(n36076), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=311, LSE_RLINE=311 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i38566_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n14011), 
         .Z(n54869)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38566_4_lut_then_3_lut.init = 16'h1010;
    CCU2D add_3134_33 (.A0(bit_counter[31]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47951), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_33.INIT0 = 16'h5999;
    defparam add_3134_33.INIT1 = 16'h0000;
    defparam add_3134_33.INJECT1_0 = "NO";
    defparam add_3134_33.INJECT1_1 = "NO";
    CCU2D add_3134_31 (.A0(bit_counter[29]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47950), .COUT(n47951), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_31.INIT0 = 16'h5999;
    defparam add_3134_31.INIT1 = 16'h5999;
    defparam add_3134_31.INJECT1_0 = "NO";
    defparam add_3134_31.INJECT1_1 = "NO";
    CCU2D add_3134_29 (.A0(bit_counter[27]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47949), .COUT(n47950), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_29.INIT0 = 16'h5999;
    defparam add_3134_29.INIT1 = 16'h5999;
    defparam add_3134_29.INJECT1_0 = "NO";
    defparam add_3134_29.INJECT1_1 = "NO";
    CCU2D add_3134_27 (.A0(bit_counter[25]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47948), .COUT(n47949), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_27.INIT0 = 16'h5999;
    defparam add_3134_27.INIT1 = 16'h5999;
    defparam add_3134_27.INJECT1_0 = "NO";
    defparam add_3134_27.INJECT1_1 = "NO";
    CCU2D add_3134_25 (.A0(bit_counter[23]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47947), .COUT(n47948), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_25.INIT0 = 16'h5999;
    defparam add_3134_25.INIT1 = 16'h5999;
    defparam add_3134_25.INJECT1_0 = "NO";
    defparam add_3134_25.INJECT1_1 = "NO";
    CCU2D add_3134_23 (.A0(bit_counter[21]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47946), .COUT(n47947), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_23.INIT0 = 16'h5999;
    defparam add_3134_23.INIT1 = 16'h5999;
    defparam add_3134_23.INJECT1_0 = "NO";
    defparam add_3134_23.INJECT1_1 = "NO";
    CCU2D add_3134_21 (.A0(bit_counter[19]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47945), .COUT(n47946), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_21.INIT0 = 16'h5999;
    defparam add_3134_21.INIT1 = 16'h5999;
    defparam add_3134_21.INJECT1_0 = "NO";
    defparam add_3134_21.INJECT1_1 = "NO";
    CCU2D add_3134_19 (.A0(bit_counter[17]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47944), .COUT(n47945), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_19.INIT0 = 16'h5999;
    defparam add_3134_19.INIT1 = 16'h5999;
    defparam add_3134_19.INJECT1_0 = "NO";
    defparam add_3134_19.INJECT1_1 = "NO";
    CCU2D add_3134_17 (.A0(bit_counter[15]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47943), .COUT(n47944), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_17.INIT0 = 16'h5999;
    defparam add_3134_17.INIT1 = 16'h5999;
    defparam add_3134_17.INJECT1_0 = "NO";
    defparam add_3134_17.INJECT1_1 = "NO";
    CCU2D add_3134_15 (.A0(bit_counter[13]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47942), .COUT(n47943), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_15.INIT0 = 16'h5999;
    defparam add_3134_15.INIT1 = 16'h5999;
    defparam add_3134_15.INJECT1_0 = "NO";
    defparam add_3134_15.INJECT1_1 = "NO";
    CCU2D add_3134_13 (.A0(bit_counter[11]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47941), .COUT(n47942), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_13.INIT0 = 16'h5999;
    defparam add_3134_13.INIT1 = 16'h5999;
    defparam add_3134_13.INJECT1_0 = "NO";
    defparam add_3134_13.INJECT1_1 = "NO";
    CCU2D add_3134_11 (.A0(bit_counter[9]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47940), .COUT(n47941), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_11.INIT0 = 16'h5999;
    defparam add_3134_11.INIT1 = 16'h5999;
    defparam add_3134_11.INJECT1_0 = "NO";
    defparam add_3134_11.INJECT1_1 = "NO";
    CCU2D add_3134_9 (.A0(bit_counter[7]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47939), .COUT(n47940), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_9.INIT0 = 16'h5999;
    defparam add_3134_9.INIT1 = 16'h5999;
    defparam add_3134_9.INJECT1_0 = "NO";
    defparam add_3134_9.INJECT1_1 = "NO";
    CCU2D add_3134_7 (.A0(bit_counter[5]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47938), .COUT(n47939), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_7.INIT0 = 16'h5999;
    defparam add_3134_7.INIT1 = 16'h5999;
    defparam add_3134_7.INJECT1_0 = "NO";
    defparam add_3134_7.INJECT1_1 = "NO";
    CCU2D add_3134_5 (.A0(bit_counter[3]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47937), .COUT(n47938), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_5.INIT0 = 16'h5999;
    defparam add_3134_5.INIT1 = 16'h5999;
    defparam add_3134_5.INJECT1_0 = "NO";
    defparam add_3134_5.INJECT1_1 = "NO";
    CCU2D add_3134_3 (.A0(bit_counter[1]), .B0(n13976), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13976), .C1(GND_net), 
          .D1(GND_net), .CIN(n47936), .COUT(n47937), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_3.INIT0 = 16'h5999;
    defparam add_3134_3.INIT1 = 16'h5999;
    defparam add_3134_3.INJECT1_0 = "NO";
    defparam add_3134_3.INJECT1_1 = "NO";
    CCU2D add_3134_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13976), .C1(GND_net), .D1(GND_net), 
          .COUT(n47936), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3134_1.INIT0 = 16'hF000;
    defparam add_3134_1.INIT1 = 16'h5999;
    defparam add_3134_1.INJECT1_0 = "NO";
    defparam add_3134_1.INJECT1_1 = "NO";
    LUT4 mux_2790_i1_4_lut (.A(n74), .B(n15105[0]), .C(n10125), .D(n52667), 
         .Z(n10126[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2790_i1_4_lut.init = 16'hcfca;
    LUT4 i2802_3_lut (.A(state[2]), .B(state[1]), .C(n14011), .Z(n10125)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2802_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42684)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i25677_1_lut_rep_760 (.A(state[2]), .Z(n54763)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25677_1_lut_rep_760.init = 16'h5555;
    LUT4 i28643_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28643_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_2_lut_rep_628 (.A(state[1]), .B(n14011), .Z(n54631)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_628.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut_adj_299 (.A(state[1]), .B(n14011), .C(n54774), 
         .D(n54638), .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_299.init = 16'hd080;
    LUT4 i28788_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28788_2_lut.init = 16'hbbbb;
    LUT4 i28787_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_901)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28787_2_lut.init = 16'hbbbb;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53175), .B(n53354), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i29431_4_lut (.A(n7204[0]), .B(n7211), .C(state[0]), .D(n54631), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29431_4_lut.init = 16'h0322;
    LUT4 i1_4_lut_adj_300 (.A(state[2]), .B(state[0]), .C(state[1]), .D(n14011), 
         .Z(n7211)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_adj_300.init = 16'ha8a0;
    LUT4 i23888_4_lut (.A(sclk_c_enable_1840), .B(n54704), .C(n10125), 
         .D(n54580), .Z(n36080)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23888_4_lut.init = 16'haaa2;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48062), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48061), .COUT(n48062), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48060), .COUT(n48061), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48059), .COUT(n48060), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48058), .COUT(n48059), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48057), .COUT(n48058), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48056), .COUT(n48057), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48055), .COUT(n48056), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48054), .COUT(n48055), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48053), .COUT(n48054), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48052), .COUT(n48053), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48051), .COUT(n48052), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48050), .COUT(n48051), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48049), .COUT(n48050), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48048), .COUT(n48049), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48047), .COUT(n48048), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48047), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48045), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48044), .COUT(n48045), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48043), .COUT(n48044), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48042), .COUT(n48043), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48042), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    PFUMX i38887 (.BLUT(n54868), .ALUT(n54869), .C0(state[1]), .Z(state_2__N_104[1]));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U27 
//

module \WS2812(48000000,"111111111")_U27  (sclk_c, \port_status[20] , ws2813_out_c_20, 
            \Q[20] , \RdAddress[20] , GND_net);
    input sclk_c;
    output \port_status[20] ;
    output ws2813_out_c_20;
    input [23:0]\Q[20] ;
    output [8:0]\RdAddress[20] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_1460;
    wire [31:0]n11194;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire n15, sclk_c_enable_177, n54746, sclk_c_enable_178, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_182;
    wire [2:0]state_2__N_104;
    
    wire n14291, n54563, n14;
    wire [31:0]n447;
    
    wire n14256, n54898, n54623, n54757, n54627, n53229, n53230;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53233, n53231, n53232, n53234, n53380, n53381, n53382, 
        n54848, n54847, n54558, n54693;
    wire [31:0]n11018;
    
    wire n80;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire sclk_c_enable_1234, n36613, sclk_c_enable_1212;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1334;
    wire [31:0]bit_counter_31__N_172;
    
    wire n54899, n37333;
    wire [8:0]n118;
    
    wire n53376, n53377, n53378, n53379, n1, n1_adj_900, n36460, 
        n36456;
    wire [31:0]n11120;
    
    wire n54900, n54626, n11193, n52727, n54754;
    wire [2:0]n6358;
    
    wire n53228, n53227, n53226, n53225, n53224, n53223, n53221, 
        n53222, n71;
    wire [6:0]n15137;
    
    wire n37343, n42636, n4, n53235, serial_N_437;
    wire [31:0]bit_counter_31__N_204;
    
    wire n74, n48929, n48928, n48927, n48926, n48925, n48924, 
        n48146, n48923, n48145, n48922, n48144, n48921, n48920, 
        n48143, n48919, n48918, n48917, n48916, n48915, n48914, 
        n48913, n48912, n48911, n48910, n48909, n48908, n48907, 
        n48906, n48905, n48904, n48903, n48902, n48901, n48900, 
        n48142, n48141, n48899, n48898, n48140, n48139, n48138, 
        n48137, n48136, n48135, n48134, n48133, n48132, n48131, 
        n48129, n6365, n48128, n48127, n48126, n47850, n47849, 
        n47848, n47847, n47846, n47845, n47844, n47843, n47842, 
        n47841, n47840, n47839, n47838, n47837, n47836, n47835;
    
    FD1P3AX delay_counter_i0_i0 (.D(n11194[0]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[8]), .C(cur_pixel[7]), 
         .D(cur_pixel[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    FD1P3AX status_77 (.D(n54746), .SP(sclk_c_enable_177), .CK(sclk_c), 
            .Q(\port_status[20] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_178), .CK(sclk_c), 
            .Q(ws2813_out_c_20)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_182), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_182), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_182), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_560_3_lut (.A(state[2]), .B(n14291), .C(state[1]), 
         .Z(n54563)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_560_3_lut.init = 16'h4040;
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n14291), .Z(sclk_c_enable_182)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i5_3_lut (.A(cur_pixel[2]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    LUT4 mux_3008_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14256), .Z(n54898)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3008_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i1_2_lut_rep_620 (.A(state[1]), .B(n14291), .Z(n54623)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_620.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[1]), .B(n14291), .C(n54757), .D(n54627), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd080;
    L6MUX21 i38027 (.D0(n53229), .D1(n53230), .SD(bit_counter[2]), .Z(n53233));
    L6MUX21 i38028 (.D0(n53231), .D1(n53232), .SD(bit_counter[2]), .Z(n53234));
    L6MUX21 i38176 (.D0(n53380), .D1(n53381), .SD(bit_counter[2]), .Z(n53382));
    LUT4 i38474_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n14291), 
         .Z(n54848)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38474_4_lut_then_3_lut.init = 16'h1010;
    LUT4 i38474_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n14256), 
         .Z(n54847)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38474_4_lut_else_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut (.A(n54558), .B(n54757), .C(n447[8]), .D(n54693), 
         .Z(n11018[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_207 (.A(n54558), .B(n54757), .C(n447[12]), 
         .D(n54693), .Z(n11018[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_207.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_208 (.A(n54558), .B(n54757), .C(n447[9]), 
         .D(n54693), .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_208.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_209 (.A(n54558), .B(n54757), .C(n447[7]), 
         .D(n54693), .Z(n11018[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_209.init = 16'hf888;
    FD1P3IX pixel_i0 (.D(\Q[20] [0]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    FD1P3IX pixel_i23 (.D(\Q[20] [23]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[20] [22]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[20] [21]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[20] [20]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    LUT4 mux_3008_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n14291), .Z(n54899)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3008_i3_4_lut_then_4_lut.init = 16'hd1f0;
    FD1P3IX pixel_i19 (.D(\Q[20] [19]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[20] [18]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[20] [17]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[20] [16]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[20] [15]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[20] [14]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[20] [13]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[20] [12]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[20] [11]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[20] [10]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[20] [9]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[20] [8]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[20] [7]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[20] [6]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[20] [5]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[20] [4]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[20] [3]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[20] [2]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[20] [1]), .SP(sclk_c_enable_1234), .CD(n36613), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n37333), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(state[2]), .B(n37333), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_210.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_211 (.A(state[2]), .B(n37333), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_211.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_212 (.A(state[2]), .B(n37333), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_212.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_213 (.A(state[2]), .B(n37333), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_213.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_214 (.A(state[2]), .B(n37333), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_214.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_215 (.A(state[2]), .B(n37333), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_215.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_216 (.A(state[2]), .B(n37333), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_216.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_217 (.A(state[2]), .B(n37333), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_217.init = 16'h1010;
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1212), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i1 (.D(n11194[1]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n11194[3]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n11194[7]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n11194[8]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n11194[9]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n11194[12]), .SP(sclk_c_enable_1460), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    PFUMX i38174 (.BLUT(n53376), .ALUT(n53377), .C0(bit_counter[1]), .Z(n53380));
    PFUMX i38175 (.BLUT(n53378), .ALUT(n53379), .C0(bit_counter[1]), .Z(n53381));
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1234), 
            .CD(n36613), .CK(sclk_c), .Q(\RdAddress[20] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1334), .CD(n36613), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_900), .SP(sclk_c_enable_1334), .CD(n36613), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1334), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 i38570_3_lut_rep_561_4_lut (.A(state[2]), .B(n14291), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_1460)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38570_3_lut_rep_561_4_lut.init = 16'hfffb;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_1460), 
            .CD(n36460), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_1460), .CD(n36460), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_1460), .CD(n36460), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n11120[4]), .SP(sclk_c_enable_1460), 
            .CD(n36456), .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54900), .SP(sclk_c_enable_1460), .CD(n36456), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=355, LSE_RLINE=355 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i24244_2_lut_4_lut (.A(n54626), .B(state[0]), .C(state[1]), .D(n11193), 
         .Z(n36456)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i24244_2_lut_4_lut.init = 16'hfd00;
    LUT4 i1_3_lut_4_lut_4_lut_adj_218 (.A(n54757), .B(state[1]), .C(n54627), 
         .D(n54626), .Z(n52727)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_218.init = 16'hce02;
    LUT4 mux_3008_i5_4_lut_4_lut (.A(state[0]), .B(n54754), .C(n447[4]), 
         .D(n54563), .Z(n11120[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_3008_i5_4_lut_4_lut.init = 16'haad0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n54754), .C(n14256), .D(n37333), 
         .Z(n6358[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfddd;
    LUT4 i37695_2_lut_rep_624 (.A(n37333), .B(n14256), .Z(n54627)) /* synthesis lut_function=(A (B)) */ ;
    defparam i37695_2_lut_rep_624.init = 16'h8888;
    LUT4 i38022_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38022_3_lut.init = 16'hcaca;
    LUT4 i38021_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38021_3_lut.init = 16'hcaca;
    LUT4 i38020_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38020_3_lut.init = 16'hcaca;
    LUT4 i38019_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38019_3_lut.init = 16'hcaca;
    LUT4 i38018_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38018_3_lut.init = 16'hcaca;
    LUT4 i38017_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38017_3_lut.init = 16'hcaca;
    PFUMX i38023 (.BLUT(n53221), .ALUT(n53222), .C0(bit_counter[1]), .Z(n53229));
    LUT4 mux_3018_i2_4_lut (.A(n71), .B(n15137[0]), .C(n11193), .D(n52727), 
         .Z(n11194[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i2_4_lut.init = 16'hcfca;
    LUT4 i38016_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38016_3_lut.init = 16'hcaca;
    LUT4 i38015_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38015_3_lut.init = 16'hcaca;
    PFUMX i38024 (.BLUT(n53223), .ALUT(n53224), .C0(bit_counter[1]), .Z(n53230));
    LUT4 mux_3018_i4_4_lut (.A(n37343), .B(n42636), .C(n11193), .D(n4), 
         .Z(n11194[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n37333), .B(n54563), .C(n447[3]), .D(n54693), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_3018_i8_4_lut (.A(n11018[7]), .B(n42636), .C(n11193), .D(n54563), 
         .Z(n11194[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i8_4_lut.init = 16'h303a;
    LUT4 mux_3018_i9_4_lut (.A(n11018[8]), .B(n42636), .C(n11193), .D(n54563), 
         .Z(n11194[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i9_4_lut.init = 16'h303a;
    LUT4 mux_3018_i10_4_lut (.A(n80), .B(n42636), .C(n11193), .D(n54563), 
         .Z(n11194[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i10_4_lut.init = 16'h303a;
    LUT4 mux_3018_i13_4_lut (.A(n11018[12]), .B(n42636), .C(n11193), .D(n54563), 
         .Z(n11194[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i13_4_lut.init = 16'h303a;
    PFUMX i38025 (.BLUT(n53225), .ALUT(n53226), .C0(bit_counter[1]), .Z(n53231));
    LUT4 i1_2_lut_rep_623 (.A(state[2]), .B(n14291), .Z(n54626)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_623.init = 16'h4444;
    PFUMX i38026 (.BLUT(n53227), .ALUT(n53228), .C0(bit_counter[1]), .Z(n53232));
    LUT4 i1_2_lut_rep_555_3_lut (.A(n37333), .B(n14256), .C(state[1]), 
         .Z(n54558)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_555_3_lut.init = 16'h0808;
    L6MUX21 i38029 (.D0(n53233), .D1(n53234), .SD(bit_counter[3]), .Z(n53235));
    LUT4 i38173_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38173_3_lut.init = 16'hcaca;
    LUT4 i38172_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38172_3_lut.init = 16'hcaca;
    LUT4 i38171_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38171_3_lut.init = 16'hcaca;
    LUT4 i38170_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38170_3_lut.init = 16'hcaca;
    LUT4 i25133_1_lut_rep_743 (.A(state[2]), .Z(n54746)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25133_1_lut_rep_743.init = 16'h5555;
    LUT4 i29946_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i29946_3_lut_3_lut.init = 16'h5151;
    LUT4 i28796_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28796_2_lut.init = 16'hbbbb;
    LUT4 i28795_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_900)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28795_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_751 (.A(state[1]), .B(state[2]), .Z(n54754)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_751.init = 16'heeee;
    LUT4 i1_2_lut_rep_690_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54693)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_690_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_219 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_219.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_220 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_220.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15137[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_221.init = 16'h7070;
    LUT4 i1_3_lut_rep_692_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1234)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_692_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n14291), 
         .Z(sclk_c_enable_178)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i30459_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42636)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i30459_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_754 (.A(state[0]), .B(state[2]), .Z(n54757)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_754.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_222 (.A(state[0]), .B(state[2]), .C(n14256), 
         .D(state[1]), .Z(n37343)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_222.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n14256), 
         .D(state[1]), .Z(sclk_c_enable_1212)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_223.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_224.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_225 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_225.init = 16'h2020;
    LUT4 i24268_4_lut (.A(sclk_c_enable_1460), .B(n54693), .C(n11193), 
         .D(n54563), .Z(n36460)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i24268_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_adj_226 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_226.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_227 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_227.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_228.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_229 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_229.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_230.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_231 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_231.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_232 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_232.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_233 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_233.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_234 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_234.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_235 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_235.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_236 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_236.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_237 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_237.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_238 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_238.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_239 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_239.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_240 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_240.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_241.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_242 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_242.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_243 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_243.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_244 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_244.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_245 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_245.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_246 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_246.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_247 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_247.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_248 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_248.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_249 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_249.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_250 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_250.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_251 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_251.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_252 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_252.init = 16'h2020;
    LUT4 i38402_2_lut_rep_755 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1334)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38402_2_lut_rep_755.init = 16'h9999;
    LUT4 i24372_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36613)) /* synthesis lut_function=(A (B)) */ ;
    defparam i24372_2_lut_2_lut.init = 16'h8888;
    CCU2D add_33930_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48929), 
          .S0(n14291));
    defparam add_33930_cout.INIT0 = 16'h0000;
    defparam add_33930_cout.INIT1 = 16'h0000;
    defparam add_33930_cout.INJECT1_0 = "NO";
    defparam add_33930_cout.INJECT1_1 = "NO";
    CCU2D add_33930_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48928), .COUT(n48929));
    defparam add_33930_31.INIT0 = 16'hf555;
    defparam add_33930_31.INIT1 = 16'h5555;
    defparam add_33930_31.INJECT1_0 = "NO";
    defparam add_33930_31.INJECT1_1 = "NO";
    CCU2D add_33930_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48927), .COUT(n48928));
    defparam add_33930_29.INIT0 = 16'hf555;
    defparam add_33930_29.INIT1 = 16'hf555;
    defparam add_33930_29.INJECT1_0 = "NO";
    defparam add_33930_29.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    CCU2D add_33930_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48926), .COUT(n48927));
    defparam add_33930_27.INIT0 = 16'hf555;
    defparam add_33930_27.INIT1 = 16'hf555;
    defparam add_33930_27.INJECT1_0 = "NO";
    defparam add_33930_27.INJECT1_1 = "NO";
    CCU2D add_33930_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48925), .COUT(n48926));
    defparam add_33930_25.INIT0 = 16'hf555;
    defparam add_33930_25.INIT1 = 16'hf555;
    defparam add_33930_25.INJECT1_0 = "NO";
    defparam add_33930_25.INJECT1_1 = "NO";
    CCU2D add_33930_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48924), .COUT(n48925));
    defparam add_33930_23.INIT0 = 16'hf555;
    defparam add_33930_23.INIT1 = 16'hf555;
    defparam add_33930_23.INJECT1_0 = "NO";
    defparam add_33930_23.INJECT1_1 = "NO";
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48146), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_33930_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48923), .COUT(n48924));
    defparam add_33930_21.INIT0 = 16'hf555;
    defparam add_33930_21.INIT1 = 16'hf555;
    defparam add_33930_21.INJECT1_0 = "NO";
    defparam add_33930_21.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48145), .COUT(n48146), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_33930_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48922), .COUT(n48923));
    defparam add_33930_19.INIT0 = 16'hf555;
    defparam add_33930_19.INIT1 = 16'hf555;
    defparam add_33930_19.INJECT1_0 = "NO";
    defparam add_33930_19.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48144), .COUT(n48145), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_33930_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48921), .COUT(n48922));
    defparam add_33930_17.INIT0 = 16'hf555;
    defparam add_33930_17.INIT1 = 16'hf555;
    defparam add_33930_17.INJECT1_0 = "NO";
    defparam add_33930_17.INJECT1_1 = "NO";
    CCU2D add_33930_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48920), .COUT(n48921));
    defparam add_33930_15.INIT0 = 16'hf555;
    defparam add_33930_15.INIT1 = 16'hf555;
    defparam add_33930_15.INJECT1_0 = "NO";
    defparam add_33930_15.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48143), .COUT(n48144), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_33930_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48919), .COUT(n48920));
    defparam add_33930_13.INIT0 = 16'hf555;
    defparam add_33930_13.INIT1 = 16'hf555;
    defparam add_33930_13.INJECT1_0 = "NO";
    defparam add_33930_13.INJECT1_1 = "NO";
    CCU2D add_33930_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48918), .COUT(n48919));
    defparam add_33930_11.INIT0 = 16'hf555;
    defparam add_33930_11.INIT1 = 16'hf555;
    defparam add_33930_11.INJECT1_0 = "NO";
    defparam add_33930_11.INJECT1_1 = "NO";
    CCU2D add_33930_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48917), .COUT(n48918));
    defparam add_33930_9.INIT0 = 16'hf555;
    defparam add_33930_9.INIT1 = 16'hf555;
    defparam add_33930_9.INJECT1_0 = "NO";
    defparam add_33930_9.INJECT1_1 = "NO";
    CCU2D add_33930_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48916), .COUT(n48917));
    defparam add_33930_7.INIT0 = 16'hf555;
    defparam add_33930_7.INIT1 = 16'hf555;
    defparam add_33930_7.INJECT1_0 = "NO";
    defparam add_33930_7.INJECT1_1 = "NO";
    CCU2D add_33930_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48915), .COUT(n48916));
    defparam add_33930_5.INIT0 = 16'hf555;
    defparam add_33930_5.INIT1 = 16'hf555;
    defparam add_33930_5.INJECT1_0 = "NO";
    defparam add_33930_5.INJECT1_1 = "NO";
    CCU2D add_33930_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48914), .COUT(n48915));
    defparam add_33930_3.INIT0 = 16'hf555;
    defparam add_33930_3.INIT1 = 16'hf555;
    defparam add_33930_3.INJECT1_0 = "NO";
    defparam add_33930_3.INJECT1_1 = "NO";
    CCU2D add_33930_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48914));
    defparam add_33930_1.INIT0 = 16'hF000;
    defparam add_33930_1.INIT1 = 16'ha666;
    defparam add_33930_1.INJECT1_0 = "NO";
    defparam add_33930_1.INJECT1_1 = "NO";
    CCU2D add_33931_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48913), 
          .S0(n14256));
    defparam add_33931_cout.INIT0 = 16'h0000;
    defparam add_33931_cout.INIT1 = 16'h0000;
    defparam add_33931_cout.INJECT1_0 = "NO";
    defparam add_33931_cout.INJECT1_1 = "NO";
    CCU2D add_33931_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48912), .COUT(n48913));
    defparam add_33931_31.INIT0 = 16'hf555;
    defparam add_33931_31.INIT1 = 16'h5555;
    defparam add_33931_31.INJECT1_0 = "NO";
    defparam add_33931_31.INJECT1_1 = "NO";
    CCU2D add_33931_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48911), .COUT(n48912));
    defparam add_33931_29.INIT0 = 16'hf555;
    defparam add_33931_29.INIT1 = 16'hf555;
    defparam add_33931_29.INJECT1_0 = "NO";
    defparam add_33931_29.INJECT1_1 = "NO";
    CCU2D add_33931_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48910), .COUT(n48911));
    defparam add_33931_27.INIT0 = 16'hf555;
    defparam add_33931_27.INIT1 = 16'hf555;
    defparam add_33931_27.INJECT1_0 = "NO";
    defparam add_33931_27.INJECT1_1 = "NO";
    CCU2D add_33931_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48909), .COUT(n48910));
    defparam add_33931_25.INIT0 = 16'hf555;
    defparam add_33931_25.INIT1 = 16'hf555;
    defparam add_33931_25.INJECT1_0 = "NO";
    defparam add_33931_25.INJECT1_1 = "NO";
    CCU2D add_33931_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48908), .COUT(n48909));
    defparam add_33931_23.INIT0 = 16'hf555;
    defparam add_33931_23.INIT1 = 16'hf555;
    defparam add_33931_23.INJECT1_0 = "NO";
    defparam add_33931_23.INJECT1_1 = "NO";
    CCU2D add_33931_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48907), .COUT(n48908));
    defparam add_33931_21.INIT0 = 16'hf555;
    defparam add_33931_21.INIT1 = 16'hf555;
    defparam add_33931_21.INJECT1_0 = "NO";
    defparam add_33931_21.INJECT1_1 = "NO";
    CCU2D add_33931_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48906), .COUT(n48907));
    defparam add_33931_19.INIT0 = 16'hf555;
    defparam add_33931_19.INIT1 = 16'hf555;
    defparam add_33931_19.INJECT1_0 = "NO";
    defparam add_33931_19.INJECT1_1 = "NO";
    CCU2D add_33931_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48905), .COUT(n48906));
    defparam add_33931_17.INIT0 = 16'hf555;
    defparam add_33931_17.INIT1 = 16'hf555;
    defparam add_33931_17.INJECT1_0 = "NO";
    defparam add_33931_17.INJECT1_1 = "NO";
    CCU2D add_33931_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48904), .COUT(n48905));
    defparam add_33931_15.INIT0 = 16'hf555;
    defparam add_33931_15.INIT1 = 16'hf555;
    defparam add_33931_15.INJECT1_0 = "NO";
    defparam add_33931_15.INJECT1_1 = "NO";
    CCU2D add_33931_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48903), .COUT(n48904));
    defparam add_33931_13.INIT0 = 16'hf555;
    defparam add_33931_13.INIT1 = 16'hf555;
    defparam add_33931_13.INJECT1_0 = "NO";
    defparam add_33931_13.INJECT1_1 = "NO";
    CCU2D add_33931_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48902), .COUT(n48903));
    defparam add_33931_11.INIT0 = 16'hf555;
    defparam add_33931_11.INIT1 = 16'hf555;
    defparam add_33931_11.INJECT1_0 = "NO";
    defparam add_33931_11.INJECT1_1 = "NO";
    CCU2D add_33931_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48901), .COUT(n48902));
    defparam add_33931_9.INIT0 = 16'hf555;
    defparam add_33931_9.INIT1 = 16'hf555;
    defparam add_33931_9.INJECT1_0 = "NO";
    defparam add_33931_9.INJECT1_1 = "NO";
    CCU2D add_33931_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48900), .COUT(n48901));
    defparam add_33931_7.INIT0 = 16'hf555;
    defparam add_33931_7.INIT1 = 16'hf555;
    defparam add_33931_7.INJECT1_0 = "NO";
    defparam add_33931_7.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48142), .COUT(n48143), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48141), .COUT(n48142), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_33931_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48899), .COUT(n48900));
    defparam add_33931_5.INIT0 = 16'hf555;
    defparam add_33931_5.INIT1 = 16'hf555;
    defparam add_33931_5.INJECT1_0 = "NO";
    defparam add_33931_5.INJECT1_1 = "NO";
    CCU2D add_33931_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48898), .COUT(n48899));
    defparam add_33931_3.INIT0 = 16'hf555;
    defparam add_33931_3.INIT1 = 16'hf555;
    defparam add_33931_3.INJECT1_0 = "NO";
    defparam add_33931_3.INJECT1_1 = "NO";
    CCU2D add_33931_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48898));
    defparam add_33931_1.INIT0 = 16'hF000;
    defparam add_33931_1.INIT1 = 16'ha666;
    defparam add_33931_1.INJECT1_0 = "NO";
    defparam add_33931_1.INJECT1_1 = "NO";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53235), .B(n53382), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48140), .COUT(n48141), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48139), .COUT(n48140), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48138), .COUT(n48139), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48137), .COUT(n48138), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48136), .COUT(n48137), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48135), .COUT(n48136), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48134), .COUT(n48135), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48133), .COUT(n48134), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48132), .COUT(n48133), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48131), .COUT(n48132), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48131), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    PFUMX i38873 (.BLUT(n54847), .ALUT(n54848), .C0(state[1]), .Z(state_2__N_104[1]));
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48129), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    LUT4 i29455_4_lut (.A(n6358[0]), .B(n6365), .C(state[0]), .D(n54623), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29455_4_lut.init = 16'h0322;
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48128), .COUT(n48129), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48127), .COUT(n48128), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48126), .COUT(n48127), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48126), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_253 (.A(state[2]), .B(state[0]), .C(state[1]), .D(n14291), 
         .Z(n6365)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_adj_253.init = 16'ha8a0;
    CCU2D add_3142_33 (.A0(bit_counter[31]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47850), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_33.INIT0 = 16'h5999;
    defparam add_3142_33.INIT1 = 16'h0000;
    defparam add_3142_33.INJECT1_0 = "NO";
    defparam add_3142_33.INJECT1_1 = "NO";
    CCU2D add_3142_31 (.A0(bit_counter[29]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47849), .COUT(n47850), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_31.INIT0 = 16'h5999;
    defparam add_3142_31.INIT1 = 16'h5999;
    defparam add_3142_31.INJECT1_0 = "NO";
    defparam add_3142_31.INJECT1_1 = "NO";
    CCU2D add_3142_29 (.A0(bit_counter[27]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47848), .COUT(n47849), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_29.INIT0 = 16'h5999;
    defparam add_3142_29.INIT1 = 16'h5999;
    defparam add_3142_29.INJECT1_0 = "NO";
    defparam add_3142_29.INJECT1_1 = "NO";
    CCU2D add_3142_27 (.A0(bit_counter[25]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47847), .COUT(n47848), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_27.INIT0 = 16'h5999;
    defparam add_3142_27.INIT1 = 16'h5999;
    defparam add_3142_27.INJECT1_0 = "NO";
    defparam add_3142_27.INJECT1_1 = "NO";
    CCU2D add_3142_25 (.A0(bit_counter[23]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47846), .COUT(n47847), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_25.INIT0 = 16'h5999;
    defparam add_3142_25.INIT1 = 16'h5999;
    defparam add_3142_25.INJECT1_0 = "NO";
    defparam add_3142_25.INJECT1_1 = "NO";
    CCU2D add_3142_23 (.A0(bit_counter[21]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47845), .COUT(n47846), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_23.INIT0 = 16'h5999;
    defparam add_3142_23.INIT1 = 16'h5999;
    defparam add_3142_23.INJECT1_0 = "NO";
    defparam add_3142_23.INJECT1_1 = "NO";
    CCU2D add_3142_21 (.A0(bit_counter[19]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47844), .COUT(n47845), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_21.INIT0 = 16'h5999;
    defparam add_3142_21.INIT1 = 16'h5999;
    defparam add_3142_21.INJECT1_0 = "NO";
    defparam add_3142_21.INJECT1_1 = "NO";
    CCU2D add_3142_19 (.A0(bit_counter[17]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47843), .COUT(n47844), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_19.INIT0 = 16'h5999;
    defparam add_3142_19.INIT1 = 16'h5999;
    defparam add_3142_19.INJECT1_0 = "NO";
    defparam add_3142_19.INJECT1_1 = "NO";
    LUT4 mux_3018_i1_4_lut (.A(n74), .B(n15137[0]), .C(n11193), .D(n52727), 
         .Z(n11194[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_3018_i1_4_lut.init = 16'hcfca;
    LUT4 i3030_3_lut (.A(state[2]), .B(state[1]), .C(n14291), .Z(n11193)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i3030_3_lut.init = 16'ha8a8;
    CCU2D add_3142_17 (.A0(bit_counter[15]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47842), .COUT(n47843), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_17.INIT0 = 16'h5999;
    defparam add_3142_17.INIT1 = 16'h5999;
    defparam add_3142_17.INJECT1_0 = "NO";
    defparam add_3142_17.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[4]), .C(n14), .D(cur_pixel[6]), 
         .Z(n37333)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    CCU2D add_3142_15 (.A0(bit_counter[13]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47841), .COUT(n47842), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_15.INIT0 = 16'h5999;
    defparam add_3142_15.INIT1 = 16'h5999;
    defparam add_3142_15.INJECT1_0 = "NO";
    defparam add_3142_15.INJECT1_1 = "NO";
    CCU2D add_3142_13 (.A0(bit_counter[11]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47840), .COUT(n47841), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_13.INIT0 = 16'h5999;
    defparam add_3142_13.INIT1 = 16'h5999;
    defparam add_3142_13.INJECT1_0 = "NO";
    defparam add_3142_13.INJECT1_1 = "NO";
    CCU2D add_3142_11 (.A0(bit_counter[9]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47839), .COUT(n47840), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_11.INIT0 = 16'h5999;
    defparam add_3142_11.INIT1 = 16'h5999;
    defparam add_3142_11.INJECT1_0 = "NO";
    defparam add_3142_11.INJECT1_1 = "NO";
    CCU2D add_3142_9 (.A0(bit_counter[7]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47838), .COUT(n47839), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_9.INIT0 = 16'h5999;
    defparam add_3142_9.INIT1 = 16'h5999;
    defparam add_3142_9.INJECT1_0 = "NO";
    defparam add_3142_9.INJECT1_1 = "NO";
    CCU2D add_3142_7 (.A0(bit_counter[5]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47837), .COUT(n47838), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_7.INIT0 = 16'h5999;
    defparam add_3142_7.INIT1 = 16'h5999;
    defparam add_3142_7.INJECT1_0 = "NO";
    defparam add_3142_7.INJECT1_1 = "NO";
    CCU2D add_3142_5 (.A0(bit_counter[3]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47836), .COUT(n47837), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_5.INIT0 = 16'h5999;
    defparam add_3142_5.INIT1 = 16'h5999;
    defparam add_3142_5.INJECT1_0 = "NO";
    defparam add_3142_5.INJECT1_1 = "NO";
    CCU2D add_3142_3 (.A0(bit_counter[1]), .B0(n14256), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n14256), .C1(GND_net), 
          .D1(GND_net), .CIN(n47835), .COUT(n47836), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_3.INIT0 = 16'h5999;
    defparam add_3142_3.INIT1 = 16'h5999;
    defparam add_3142_3.INJECT1_0 = "NO";
    defparam add_3142_3.INJECT1_1 = "NO";
    CCU2D add_3142_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n14256), .C1(GND_net), .D1(GND_net), 
          .COUT(n47835), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3142_1.INIT0 = 16'hF000;
    defparam add_3142_1.INIT1 = 16'h5999;
    defparam add_3142_1.INJECT1_0 = "NO";
    defparam add_3142_1.INJECT1_1 = "NO";
    PFUMX i38907 (.BLUT(n54898), .ALUT(n54899), .C0(state[1]), .Z(n54900));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U34 
//

module \WS2812(48000000,"111111111")_U34  (GND_net, sclk_c, \port_status[14] , 
            ws2813_out_c_14, \Q[14] , \RdAddress[14] );
    input GND_net;
    input sclk_c;
    output \port_status[14] ;
    output ws2813_out_c_14;
    input [23:0]\Q[14] ;
    output [8:0]\RdAddress[14] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n48017;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    wire [31:0]n447;
    
    wire n48018, n48016, sclk_c_enable_2030;
    wire [31:0]n9592;
    
    wire sclk_c_enable_130, n54772, sclk_c_enable_131, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_135;
    wire [2:0]state_2__N_104;
    
    wire n48015, n48014, n48013, n48012, n48011, n48010, n48009, 
        n48008, n54707, n13871, n7755, n48007, sclk_c_enable_1848, 
        n69, n48006, n53139, n53140;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53143, n48005, n68, n53141, n53142, n53144, n36068, 
        n54783, n13836, n38153, sclk_c_enable_1815;
    wire [31:0]bit_counter_31__N_204;
    wire [31:0]bit_counter_31__N_172;
    
    wire n48003;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]n118;
    
    wire n54643, n54588, n42580, n54644, n54578, n103, n54959, 
        n54958;
    wire [31:0]n9416;
    
    wire n76, serial_N_437, n53338, n53339, n53340, n48002;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_1879, n48001, n48000, n54703, n54853, n54854, 
        n54855, n53131, n53132, n53133, n53134, n53135, n53136, 
        n53137, n53138, n9591, n35890, n53337, n53336, n53335, 
        n53334, n52658, n35886, n47983, n47982, n47981, n47980, 
        n47979, n47978, n47977, n53145, n47976, n47975, n47974, 
        n47973, n47972, n47971, n47970, n47969, n47968, n36039, 
        n49023, n49022, n49021, n49020, n49019, n49018, n49017, 
        n49016, n49015, n1, n49014, n1_adj_899, n49013, n49012, 
        n49011, n49010, n49009;
    wire [6:0]n15089;
    
    wire n49008, n15, n14, n54960, n4, n48945, n48944, n48943, 
        n48942, n48941, n48940, n48939, n48938, n48937, n48936, 
        n48935, n48934, n48933, n48932, n48931, n48930, n48020, 
        n48019;
    
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48017), .COUT(n48018), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48016), .COUT(n48017), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    FD1P3AX delay_counter_i0_i0 (.D(n9592[0]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54772), .SP(sclk_c_enable_130), .CK(sclk_c), 
            .Q(\port_status[14] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_131), .CK(sclk_c), 
            .Q(ws2813_out_c_14)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_135), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_135), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_135), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48015), .COUT(n48016), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48014), .COUT(n48015), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48013), .COUT(n48014), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48012), .COUT(n48013), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48011), .COUT(n48012), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48010), .COUT(n48011), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48009), .COUT(n48010), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48008), .COUT(n48009), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_704_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54707)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_704_3_lut.init = 16'hefef;
    LUT4 i1_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(n13871), .Z(n7755)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hec88;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n13871), 
         .Z(sclk_c_enable_131)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48007), .COUT(n48008), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_683_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_1848)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_683_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n69)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48006), .COUT(n48007), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    L6MUX21 i37937 (.D0(n53139), .D1(n53140), .SD(bit_counter[2]), .Z(n53143));
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48005), .COUT(n48006), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_164 (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n68)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_164.init = 16'he0f0;
    L6MUX21 i37938 (.D0(n53141), .D1(n53142), .SD(bit_counter[2]), .Z(n53144));
    LUT4 i38449_3_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13871), .Z(sclk_c_enable_135)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38449_3_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i23919_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n36068)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i23919_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_780 (.A(state[0]), .B(state[2]), .Z(n54783)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_780.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_165 (.A(state[0]), .B(state[2]), .C(n13836), 
         .D(state[1]), .Z(n38153)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut_adj_165.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13836), 
         .D(state[1]), .Z(sclk_c_enable_1815)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_166 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_166.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_167 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_167.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_168 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_168.init = 16'h2020;
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48005), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_169 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_169.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_170 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_170.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_171 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_171.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_172 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_172.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_173 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_173.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_174 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_174.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_175 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_175.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_176 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_176.init = 16'h2020;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48003), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_177 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_177.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_178 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_178.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_179 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_179.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_180 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_180.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_181 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_181.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_182 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_182.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_183 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_183.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_184 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_184.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_185 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_185.init = 16'h2020;
    LUT4 i1_2_lut_rep_640 (.A(state[2]), .B(n13871), .Z(n54643)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_640.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_adj_186 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_186.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_187 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_187.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_188 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_188.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_189 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_189.init = 16'h2020;
    LUT4 i1_2_lut_rep_585_3_lut (.A(state[2]), .B(n13871), .C(state[1]), 
         .Z(n54588)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_585_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_190 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_190.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_191 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_191.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_192 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_192.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_193 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_193.init = 16'h2020;
    LUT4 i38585_3_lut_rep_586_4_lut (.A(state[2]), .B(n13871), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2030)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38585_3_lut_rep_586_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_adj_194 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_194.init = 16'h2020;
    LUT4 i1_2_lut_rep_641 (.A(n42580), .B(n13836), .Z(n54644)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_641.init = 16'h8888;
    LUT4 i1_2_lut_rep_575_3_lut (.A(n42580), .B(n13836), .C(state[1]), 
         .Z(n54578)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_575_3_lut.init = 16'h0808;
    LUT4 i107_3_lut_4_lut (.A(n42580), .B(n13836), .C(n54707), .D(n447[12]), 
         .Z(n103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i107_3_lut_4_lut.init = 16'hf808;
    LUT4 i25952_1_lut_rep_769 (.A(state[2]), .Z(n54772)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i25952_1_lut_rep_769.init = 16'h5555;
    LUT4 mux_2666_i5_4_lut_4_lut_then_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13871), .Z(n54959)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2666_i5_4_lut_4_lut_then_4_lut.init = 16'he4e0;
    LUT4 mux_2666_i5_4_lut_4_lut_else_4_lut (.A(state[2]), .B(state[1]), 
         .C(n447[4]), .D(n13871), .Z(n54958)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2666_i5_4_lut_4_lut_else_4_lut.init = 16'hb0f0;
    LUT4 i1_3_lut_4_lut (.A(n54578), .B(n54783), .C(n447[7]), .D(n54707), 
         .Z(n9416[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_195 (.A(n54578), .B(n54783), .C(n447[8]), 
         .D(n54707), .Z(n9416[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_195.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_196 (.A(n54578), .B(n54783), .C(n447[9]), 
         .D(n54707), .Z(n76)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_196.init = 16'hf888;
    LUT4 i28664_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28664_3_lut_3_lut.init = 16'h5151;
    L6MUX21 i38134 (.D0(n53338), .D1(n53339), .SD(bit_counter[2]), .Z(n53340));
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48002), .COUT(n48003), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    FD1P3AX delay_counter_i0_i1 (.D(n9592[1]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n9592[3]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n9592[7]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n9592[8]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n9592[9]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n9592[12]), .SP(sclk_c_enable_2030), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3IX pixel_i0 (.D(\Q[14] [0]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_197 (.A(state[2]), .B(n42580), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_197.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_198 (.A(state[2]), .B(n42580), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_198.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_199 (.A(state[2]), .B(n42580), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_199.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_200 (.A(state[2]), .B(n42580), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_200.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_201 (.A(state[2]), .B(n42580), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_201.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_202 (.A(state[2]), .B(n42580), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_202.init = 16'h1010;
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48001), .COUT(n48002), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_203 (.A(state[2]), .B(n42580), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_203.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_204 (.A(state[2]), .B(n42580), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_204.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_205 (.A(state[2]), .B(n42580), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_205.init = 16'h1010;
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48000), .COUT(n48001), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    LUT4 mux_2281_i2_4_lut_4_lut (.A(n54703), .B(n54707), .C(n7755), .D(n13836), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2281_i2_4_lut_4_lut.init = 16'h5053;
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n48000), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    PFUMX i38877 (.BLUT(n54853), .ALUT(n54854), .C0(state[1]), .Z(n54855));
    PFUMX i37933 (.BLUT(n53131), .ALUT(n53132), .C0(bit_counter[1]), .Z(n53139));
    PFUMX i37934 (.BLUT(n53133), .ALUT(n53134), .C0(bit_counter[1]), .Z(n53140));
    PFUMX i37935 (.BLUT(n53135), .ALUT(n53136), .C0(bit_counter[1]), .Z(n53141));
    PFUMX i37936 (.BLUT(n53137), .ALUT(n53138), .C0(bit_counter[1]), .Z(n53142));
    LUT4 i23698_4_lut (.A(sclk_c_enable_2030), .B(n54707), .C(n9591), 
         .D(n54588), .Z(n35890)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23698_4_lut.init = 16'haaa2;
    LUT4 mux_2666_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13871), .Z(n54854)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2666_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2666_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13836), .Z(n54853)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2666_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i38131_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38131_3_lut.init = 16'hcaca;
    LUT4 i38130_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38130_3_lut.init = 16'hcaca;
    LUT4 i38129_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38129_3_lut.init = 16'hcaca;
    LUT4 i38128_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38128_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n54783), .B(state[1]), .C(n54644), .D(n54643), 
         .Z(n52658)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hce02;
    LUT4 i23674_2_lut_4_lut (.A(n54643), .B(state[0]), .C(state[1]), .D(n9591), 
         .Z(n35886)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23674_2_lut_4_lut.init = 16'hfd00;
    CCU2D add_3130_33 (.A0(bit_counter[31]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47983), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_33.INIT0 = 16'h5999;
    defparam add_3130_33.INIT1 = 16'h0000;
    defparam add_3130_33.INJECT1_0 = "NO";
    defparam add_3130_33.INJECT1_1 = "NO";
    LUT4 i37932_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37932_3_lut.init = 16'hcaca;
    LUT4 i37931_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37931_3_lut.init = 16'hcaca;
    LUT4 i37930_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37930_3_lut.init = 16'hcaca;
    LUT4 i37929_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37929_3_lut.init = 16'hcaca;
    LUT4 i37928_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37928_3_lut.init = 16'hcaca;
    LUT4 i37927_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37927_3_lut.init = 16'hcaca;
    LUT4 i37926_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37926_3_lut.init = 16'hcaca;
    LUT4 i37925_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37925_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(state[1]), .B(n54644), .C(n13871), .D(n54783), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut_4_lut.init = 16'he400;
    CCU2D add_3130_31 (.A0(bit_counter[29]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47982), .COUT(n47983), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_31.INIT0 = 16'h5999;
    defparam add_3130_31.INIT1 = 16'h5999;
    defparam add_3130_31.INJECT1_0 = "NO";
    defparam add_3130_31.INJECT1_1 = "NO";
    CCU2D add_3130_29 (.A0(bit_counter[27]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47981), .COUT(n47982), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_29.INIT0 = 16'h5999;
    defparam add_3130_29.INIT1 = 16'h5999;
    defparam add_3130_29.INJECT1_0 = "NO";
    defparam add_3130_29.INJECT1_1 = "NO";
    CCU2D add_3130_27 (.A0(bit_counter[25]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47980), .COUT(n47981), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_27.INIT0 = 16'h5999;
    defparam add_3130_27.INIT1 = 16'h5999;
    defparam add_3130_27.INJECT1_0 = "NO";
    defparam add_3130_27.INJECT1_1 = "NO";
    CCU2D add_3130_25 (.A0(bit_counter[23]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47979), .COUT(n47980), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_25.INIT0 = 16'h5999;
    defparam add_3130_25.INIT1 = 16'h5999;
    defparam add_3130_25.INJECT1_0 = "NO";
    defparam add_3130_25.INJECT1_1 = "NO";
    CCU2D add_3130_23 (.A0(bit_counter[21]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47978), .COUT(n47979), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_23.INIT0 = 16'h5999;
    defparam add_3130_23.INIT1 = 16'h5999;
    defparam add_3130_23.INJECT1_0 = "NO";
    defparam add_3130_23.INJECT1_1 = "NO";
    CCU2D add_3130_21 (.A0(bit_counter[19]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47977), .COUT(n47978), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_21.INIT0 = 16'h5999;
    defparam add_3130_21.INIT1 = 16'h5999;
    defparam add_3130_21.INJECT1_0 = "NO";
    defparam add_3130_21.INJECT1_1 = "NO";
    L6MUX21 i37939 (.D0(n53143), .D1(n53144), .SD(bit_counter[3]), .Z(n53145));
    CCU2D add_3130_19 (.A0(bit_counter[17]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47976), .COUT(n47977), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_19.INIT0 = 16'h5999;
    defparam add_3130_19.INIT1 = 16'h5999;
    defparam add_3130_19.INJECT1_0 = "NO";
    defparam add_3130_19.INJECT1_1 = "NO";
    CCU2D add_3130_17 (.A0(bit_counter[15]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47975), .COUT(n47976), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_17.INIT0 = 16'h5999;
    defparam add_3130_17.INIT1 = 16'h5999;
    defparam add_3130_17.INJECT1_0 = "NO";
    defparam add_3130_17.INJECT1_1 = "NO";
    CCU2D add_3130_15 (.A0(bit_counter[13]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47974), .COUT(n47975), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_15.INIT0 = 16'h5999;
    defparam add_3130_15.INIT1 = 16'h5999;
    defparam add_3130_15.INJECT1_0 = "NO";
    defparam add_3130_15.INJECT1_1 = "NO";
    CCU2D add_3130_13 (.A0(bit_counter[11]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47973), .COUT(n47974), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_13.INIT0 = 16'h5999;
    defparam add_3130_13.INIT1 = 16'h5999;
    defparam add_3130_13.INJECT1_0 = "NO";
    defparam add_3130_13.INJECT1_1 = "NO";
    CCU2D add_3130_11 (.A0(bit_counter[9]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47972), .COUT(n47973), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_11.INIT0 = 16'h5999;
    defparam add_3130_11.INIT1 = 16'h5999;
    defparam add_3130_11.INJECT1_0 = "NO";
    defparam add_3130_11.INJECT1_1 = "NO";
    CCU2D add_3130_9 (.A0(bit_counter[7]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47971), .COUT(n47972), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_9.INIT0 = 16'h5999;
    defparam add_3130_9.INIT1 = 16'h5999;
    defparam add_3130_9.INJECT1_0 = "NO";
    defparam add_3130_9.INJECT1_1 = "NO";
    PFUMX i38132 (.BLUT(n53334), .ALUT(n53335), .C0(bit_counter[1]), .Z(n53338));
    PFUMX i38133 (.BLUT(n53336), .ALUT(n53337), .C0(bit_counter[1]), .Z(n53339));
    CCU2D add_3130_7 (.A0(bit_counter[5]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47970), .COUT(n47971), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_7.INIT0 = 16'h5999;
    defparam add_3130_7.INIT1 = 16'h5999;
    defparam add_3130_7.INJECT1_0 = "NO";
    defparam add_3130_7.INJECT1_1 = "NO";
    CCU2D add_3130_5 (.A0(bit_counter[3]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47969), .COUT(n47970), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_5.INIT0 = 16'h5999;
    defparam add_3130_5.INIT1 = 16'h5999;
    defparam add_3130_5.INJECT1_0 = "NO";
    defparam add_3130_5.INJECT1_1 = "NO";
    CCU2D add_3130_3 (.A0(bit_counter[1]), .B0(n13836), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13836), .C1(GND_net), 
          .D1(GND_net), .CIN(n47968), .COUT(n47969), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_3.INIT0 = 16'h5999;
    defparam add_3130_3.INIT1 = 16'h5999;
    defparam add_3130_3.INJECT1_0 = "NO";
    defparam add_3130_3.INJECT1_1 = "NO";
    CCU2D add_3130_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13836), .C1(GND_net), .D1(GND_net), 
          .COUT(n47968), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3130_1.INIT0 = 16'hF000;
    defparam add_3130_1.INIT1 = 16'h5999;
    defparam add_3130_1.INJECT1_0 = "NO";
    defparam add_3130_1.INJECT1_1 = "NO";
    LUT4 i38414_2_lut_rep_741 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1879)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38414_2_lut_rep_741.init = 16'h9999;
    LUT4 i23827_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n36039)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23827_2_lut_2_lut.init = 16'h8888;
    FD1P3IX pixel_i23 (.D(\Q[14] [23]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[14] [22]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[14] [21]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[14] [20]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[14] [19]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[14] [18]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[14] [17]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[14] [16]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[14] [15]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[14] [14]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[14] [13]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[14] [12]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[14] [11]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[14] [10]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[14] [9]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[14] [8]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[14] [7]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[14] [6]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[14] [5]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[14] [4]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[14] [3]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[14] [2]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[14] [1]), .SP(sclk_c_enable_1848), .CD(n36068), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1815), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1848), 
            .CD(n36068), .CK(sclk_c), .Q(\RdAddress[14] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_700_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54703)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_rep_700_3_lut.init = 16'hf8f8;
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    CCU2D add_33902_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49023), 
          .S0(n13871));
    defparam add_33902_cout.INIT0 = 16'h0000;
    defparam add_33902_cout.INIT1 = 16'h0000;
    defparam add_33902_cout.INJECT1_0 = "NO";
    defparam add_33902_cout.INJECT1_1 = "NO";
    CCU2D add_33902_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49022), .COUT(n49023));
    defparam add_33902_31.INIT0 = 16'hf555;
    defparam add_33902_31.INIT1 = 16'h5555;
    defparam add_33902_31.INJECT1_0 = "NO";
    defparam add_33902_31.INJECT1_1 = "NO";
    CCU2D add_33902_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49021), .COUT(n49022));
    defparam add_33902_29.INIT0 = 16'hf555;
    defparam add_33902_29.INIT1 = 16'hf555;
    defparam add_33902_29.INJECT1_0 = "NO";
    defparam add_33902_29.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    CCU2D add_33902_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49020), .COUT(n49021));
    defparam add_33902_27.INIT0 = 16'hf555;
    defparam add_33902_27.INIT1 = 16'hf555;
    defparam add_33902_27.INJECT1_0 = "NO";
    defparam add_33902_27.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    CCU2D add_33902_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49019), .COUT(n49020));
    defparam add_33902_25.INIT0 = 16'hf555;
    defparam add_33902_25.INIT1 = 16'hf555;
    defparam add_33902_25.INJECT1_0 = "NO";
    defparam add_33902_25.INJECT1_1 = "NO";
    CCU2D add_33902_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49018), .COUT(n49019));
    defparam add_33902_23.INIT0 = 16'hf555;
    defparam add_33902_23.INIT1 = 16'hf555;
    defparam add_33902_23.INJECT1_0 = "NO";
    defparam add_33902_23.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    CCU2D add_33902_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49017), .COUT(n49018));
    defparam add_33902_21.INIT0 = 16'hf555;
    defparam add_33902_21.INIT1 = 16'hf555;
    defparam add_33902_21.INJECT1_0 = "NO";
    defparam add_33902_21.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    CCU2D add_33902_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49016), .COUT(n49017));
    defparam add_33902_19.INIT0 = 16'hf555;
    defparam add_33902_19.INIT1 = 16'hf555;
    defparam add_33902_19.INJECT1_0 = "NO";
    defparam add_33902_19.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    CCU2D add_33902_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49015), .COUT(n49016));
    defparam add_33902_17.INIT0 = 16'hf555;
    defparam add_33902_17.INIT1 = 16'hf555;
    defparam add_33902_17.INJECT1_0 = "NO";
    defparam add_33902_17.INJECT1_1 = "NO";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1879), .CD(n36039), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    CCU2D add_33902_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49014), .COUT(n49015));
    defparam add_33902_15.INIT0 = 16'hf555;
    defparam add_33902_15.INIT1 = 16'hf555;
    defparam add_33902_15.INJECT1_0 = "NO";
    defparam add_33902_15.INJECT1_1 = "NO";
    FD1P3IX bit_counter_i3 (.D(n1_adj_899), .SP(sclk_c_enable_1879), .CD(n36039), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    CCU2D add_33902_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49013), .COUT(n49014));
    defparam add_33902_13.INIT0 = 16'hf555;
    defparam add_33902_13.INIT1 = 16'hf555;
    defparam add_33902_13.INJECT1_0 = "NO";
    defparam add_33902_13.INJECT1_1 = "NO";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1879), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    CCU2D add_33902_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49012), .COUT(n49013));
    defparam add_33902_11.INIT0 = 16'hf555;
    defparam add_33902_11.INIT1 = 16'hf555;
    defparam add_33902_11.INJECT1_0 = "NO";
    defparam add_33902_11.INJECT1_1 = "NO";
    CCU2D add_33902_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49011), .COUT(n49012));
    defparam add_33902_9.INIT0 = 16'hf555;
    defparam add_33902_9.INIT1 = 16'hf555;
    defparam add_33902_9.INJECT1_0 = "NO";
    defparam add_33902_9.INJECT1_1 = "NO";
    CCU2D add_33902_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49010), .COUT(n49011));
    defparam add_33902_7.INIT0 = 16'hf555;
    defparam add_33902_7.INIT1 = 16'hf555;
    defparam add_33902_7.INJECT1_0 = "NO";
    defparam add_33902_7.INJECT1_1 = "NO";
    CCU2D add_33902_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49009), .COUT(n49010));
    defparam add_33902_5.INIT0 = 16'hf555;
    defparam add_33902_5.INIT1 = 16'hf555;
    defparam add_33902_5.INJECT1_0 = "NO";
    defparam add_33902_5.INJECT1_1 = "NO";
    LUT4 mux_2676_i2_4_lut (.A(n68), .B(n15089[0]), .C(n9591), .D(n52658), 
         .Z(n9592[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i2_4_lut.init = 16'hcfca;
    CCU2D add_33902_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49008), .COUT(n49009));
    defparam add_33902_3.INIT0 = 16'hf555;
    defparam add_33902_3.INIT1 = 16'hf555;
    defparam add_33902_3.INJECT1_0 = "NO";
    defparam add_33902_3.INJECT1_1 = "NO";
    CCU2D add_33902_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n49008));
    defparam add_33902_1.INIT0 = 16'hF000;
    defparam add_33902_1.INIT1 = 16'ha666;
    defparam add_33902_1.INJECT1_0 = "NO";
    defparam add_33902_1.INJECT1_1 = "NO";
    LUT4 mux_2676_i1_4_lut (.A(n69), .B(n15089[0]), .C(n9591), .D(n52658), 
         .Z(n9592[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i1_4_lut.init = 16'hcfca;
    LUT4 i2688_3_lut (.A(state[2]), .B(state[1]), .C(n13871), .Z(n9591)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2688_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[3]), .C(n14), .D(cur_pixel[6]), 
         .Z(n42580)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[4]), .C(cur_pixel[2]), 
         .D(cur_pixel[8]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    LUT4 i5_3_lut (.A(cur_pixel[7]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2030), 
            .CD(n35890), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2030), .CD(n35890), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2030), .CD(n35890), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54960), .SP(sclk_c_enable_2030), .CD(n35886), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    LUT4 mux_2676_i4_4_lut (.A(n38153), .B(n54703), .C(n9591), .D(n4), 
         .Z(n9592[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i4_4_lut.init = 16'h3f3a;
    FD1P3IX delay_counter_i0_i2 (.D(n54855), .SP(sclk_c_enable_2030), .CD(n35886), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=289, LSE_RLINE=289 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n42580), .B(n54588), .C(n447[3]), .D(n54707), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2676_i8_4_lut (.A(n9416[7]), .B(n54703), .C(n9591), .D(n54588), 
         .Z(n9592[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i8_4_lut.init = 16'h303a;
    CCU2D add_33903_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48945), 
          .S0(n13836));
    defparam add_33903_cout.INIT0 = 16'h0000;
    defparam add_33903_cout.INIT1 = 16'h0000;
    defparam add_33903_cout.INJECT1_0 = "NO";
    defparam add_33903_cout.INJECT1_1 = "NO";
    CCU2D add_33903_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48944), .COUT(n48945));
    defparam add_33903_31.INIT0 = 16'hf555;
    defparam add_33903_31.INIT1 = 16'h5555;
    defparam add_33903_31.INJECT1_0 = "NO";
    defparam add_33903_31.INJECT1_1 = "NO";
    CCU2D add_33903_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48943), .COUT(n48944));
    defparam add_33903_29.INIT0 = 16'hf555;
    defparam add_33903_29.INIT1 = 16'hf555;
    defparam add_33903_29.INJECT1_0 = "NO";
    defparam add_33903_29.INJECT1_1 = "NO";
    CCU2D add_33903_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48942), .COUT(n48943));
    defparam add_33903_27.INIT0 = 16'hf555;
    defparam add_33903_27.INIT1 = 16'hf555;
    defparam add_33903_27.INJECT1_0 = "NO";
    defparam add_33903_27.INJECT1_1 = "NO";
    CCU2D add_33903_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48941), .COUT(n48942));
    defparam add_33903_25.INIT0 = 16'hf555;
    defparam add_33903_25.INIT1 = 16'hf555;
    defparam add_33903_25.INJECT1_0 = "NO";
    defparam add_33903_25.INJECT1_1 = "NO";
    CCU2D add_33903_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48940), .COUT(n48941));
    defparam add_33903_23.INIT0 = 16'hf555;
    defparam add_33903_23.INIT1 = 16'hf555;
    defparam add_33903_23.INJECT1_0 = "NO";
    defparam add_33903_23.INJECT1_1 = "NO";
    CCU2D add_33903_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48939), .COUT(n48940));
    defparam add_33903_21.INIT0 = 16'hf555;
    defparam add_33903_21.INIT1 = 16'hf555;
    defparam add_33903_21.INJECT1_0 = "NO";
    defparam add_33903_21.INJECT1_1 = "NO";
    CCU2D add_33903_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48938), .COUT(n48939));
    defparam add_33903_19.INIT0 = 16'hf555;
    defparam add_33903_19.INIT1 = 16'hf555;
    defparam add_33903_19.INJECT1_0 = "NO";
    defparam add_33903_19.INJECT1_1 = "NO";
    CCU2D add_33903_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48937), .COUT(n48938));
    defparam add_33903_17.INIT0 = 16'hf555;
    defparam add_33903_17.INIT1 = 16'hf555;
    defparam add_33903_17.INJECT1_0 = "NO";
    defparam add_33903_17.INJECT1_1 = "NO";
    CCU2D add_33903_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48936), .COUT(n48937));
    defparam add_33903_15.INIT0 = 16'hf555;
    defparam add_33903_15.INIT1 = 16'hf555;
    defparam add_33903_15.INJECT1_0 = "NO";
    defparam add_33903_15.INJECT1_1 = "NO";
    CCU2D add_33903_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48935), .COUT(n48936));
    defparam add_33903_13.INIT0 = 16'hf555;
    defparam add_33903_13.INIT1 = 16'hf555;
    defparam add_33903_13.INJECT1_0 = "NO";
    defparam add_33903_13.INJECT1_1 = "NO";
    CCU2D add_33903_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48934), .COUT(n48935));
    defparam add_33903_11.INIT0 = 16'hf555;
    defparam add_33903_11.INIT1 = 16'hf555;
    defparam add_33903_11.INJECT1_0 = "NO";
    defparam add_33903_11.INJECT1_1 = "NO";
    CCU2D add_33903_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48933), .COUT(n48934));
    defparam add_33903_9.INIT0 = 16'hf555;
    defparam add_33903_9.INIT1 = 16'hf555;
    defparam add_33903_9.INJECT1_0 = "NO";
    defparam add_33903_9.INJECT1_1 = "NO";
    CCU2D add_33903_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48932), .COUT(n48933));
    defparam add_33903_7.INIT0 = 16'hf555;
    defparam add_33903_7.INIT1 = 16'hf555;
    defparam add_33903_7.INJECT1_0 = "NO";
    defparam add_33903_7.INJECT1_1 = "NO";
    CCU2D add_33903_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48931), .COUT(n48932));
    defparam add_33903_5.INIT0 = 16'hf555;
    defparam add_33903_5.INIT1 = 16'hf555;
    defparam add_33903_5.INJECT1_0 = "NO";
    defparam add_33903_5.INJECT1_1 = "NO";
    CCU2D add_33903_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48930), .COUT(n48931));
    defparam add_33903_3.INIT0 = 16'hf555;
    defparam add_33903_3.INIT1 = 16'hf555;
    defparam add_33903_3.INJECT1_0 = "NO";
    defparam add_33903_3.INJECT1_1 = "NO";
    CCU2D add_33903_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48930));
    defparam add_33903_1.INIT0 = 16'hF000;
    defparam add_33903_1.INIT1 = 16'ha666;
    defparam add_33903_1.INJECT1_0 = "NO";
    defparam add_33903_1.INJECT1_1 = "NO";
    LUT4 mux_2676_i9_4_lut (.A(n9416[8]), .B(n54703), .C(n9591), .D(n54588), 
         .Z(n9592[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i9_4_lut.init = 16'h303a;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53145), .B(n53340), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2281_i1_4_lut (.A(n54644), .B(n54703), .C(n7755), .D(n54707), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2281_i1_4_lut.init = 16'h3f3a;
    LUT4 mux_2676_i10_4_lut (.A(n76), .B(n54703), .C(n9591), .D(n54588), 
         .Z(n9592[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i10_4_lut.init = 16'h303a;
    LUT4 mux_2676_i13_4_lut (.A(n54588), .B(n54703), .C(n9591), .D(n103), 
         .Z(n9592[12])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2676_i13_4_lut.init = 16'h3530;
    LUT4 i1_2_lut_3_lut_adj_206 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15089[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_206.init = 16'h7070;
    LUT4 i28784_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28784_2_lut.init = 16'hbbbb;
    LUT4 i28783_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_899)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28783_2_lut.init = 16'hbbbb;
    PFUMX i38947 (.BLUT(n54958), .ALUT(n54959), .C0(state[0]), .Z(n54960));
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48020), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48019), .COUT(n48020), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48018), .COUT(n48019), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U37 
//

module \WS2812(48000000,"111111111")_U37  (GND_net, sclk_c, \port_status[11] , 
            ws2813_out_c_11, state, n54591, \Q[11] , \RdAddress[11] );
    input GND_net;
    input sclk_c;
    output \port_status[11] ;
    output ws2813_out_c_11;
    output [2:0]state;
    input n54591;
    input [23:0]\Q[11] ;
    output [8:0]\RdAddress[11] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n48587;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire n48588, n48586, n48585, sclk_c_enable_2315;
    wire [31:0]n8746;
    
    wire n48584, sclk_c_enable_105, n54786, sclk_c_enable_106, serial_N_433, 
        sclk_c_enable_110;
    wire [2:0]state_2__N_104;
    
    wire n48583, n48582, n47804;
    wire [31:0]n447;
    
    wire n47805, n48581, n48580, n54895, n54896, n48579, n47803, 
        n47802, n48578, n53094, n53095;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53098, n53096, n53097, n53099, n47801, n47800, n47799, 
        n47798, n13661, n47796;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]n118;
    
    wire n47795, n47794, n8556, n47793, n55533, n54929, serial_N_437, 
        n54928, n54935, n54934, n13626, n11, n55538;
    wire [31:0]bit_counter_31__N_204;
    
    wire n1, n1_adj_898, n54993, n54992, n54600, n54717;
    wire [31:0]n8570;
    
    wire n42570;
    wire [6:0]n15065;
    
    wire n45, sclk_c_enable_2133, n53, n55532, sclk_c_enable_2100, 
        n38570, n53317, n53318, n53319;
    wire [31:0]bit_counter_31__N_172;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n35783;
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_2164, n8745, n35605, n53086, n53087, n53088, 
        n53089, n53090, n53091, n53092, n53093, n53316, n53315, 
        n53314, n53313, n52739, n15, n14, n53100, n48226, n48497, 
        n48225, n48496, n48224, n48495, n48223, n48494, n48222, 
        n48493, n48492, n48221, n48220, n48219, n48218, n48491, 
        n48490, n48489, n48488, n48487, n48217, n48216, n48215, 
        n48214, n48213, n48212, n48211, n48486, n48485, n48484, 
        n48483, n48482, n54936, n54994, n4, n54930, n47813, n47812, 
        n47811, n48593, n48592, n47810, n47809, n47808, n48591, 
        n47807, n48590, n47806, n48589;
    
    CCU2D add_33910_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48587), .COUT(n48588));
    defparam add_33910_21.INIT0 = 16'hf555;
    defparam add_33910_21.INIT1 = 16'hf555;
    defparam add_33910_21.INJECT1_0 = "NO";
    defparam add_33910_21.INJECT1_1 = "NO";
    CCU2D add_33910_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48586), .COUT(n48587));
    defparam add_33910_19.INIT0 = 16'hf555;
    defparam add_33910_19.INIT1 = 16'hf555;
    defparam add_33910_19.INJECT1_0 = "NO";
    defparam add_33910_19.INJECT1_1 = "NO";
    CCU2D add_33910_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48585), .COUT(n48586));
    defparam add_33910_17.INIT0 = 16'hf555;
    defparam add_33910_17.INIT1 = 16'hf555;
    defparam add_33910_17.INJECT1_0 = "NO";
    defparam add_33910_17.INJECT1_1 = "NO";
    FD1P3AX delay_counter_i0_i0 (.D(n8746[0]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    CCU2D add_33910_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48584), .COUT(n48585));
    defparam add_33910_15.INIT0 = 16'hf555;
    defparam add_33910_15.INIT1 = 16'hf555;
    defparam add_33910_15.INJECT1_0 = "NO";
    defparam add_33910_15.INJECT1_1 = "NO";
    FD1P3AX status_77 (.D(n54786), .SP(sclk_c_enable_105), .CK(sclk_c), 
            .Q(\port_status[11] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_106), .CK(sclk_c), 
            .Q(ws2813_out_c_11)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_110), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_110), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_110), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    CCU2D add_33910_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48583), .COUT(n48584));
    defparam add_33910_13.INIT0 = 16'hf555;
    defparam add_33910_13.INIT1 = 16'hf555;
    defparam add_33910_13.INJECT1_0 = "NO";
    defparam add_33910_13.INJECT1_1 = "NO";
    CCU2D add_33910_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48582), .COUT(n48583));
    defparam add_33910_11.INIT0 = 16'hf555;
    defparam add_33910_11.INIT1 = 16'hf555;
    defparam add_33910_11.INJECT1_0 = "NO";
    defparam add_33910_11.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47804), .COUT(n47805), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_33910_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48581), .COUT(n48582));
    defparam add_33910_9.INIT0 = 16'hf555;
    defparam add_33910_9.INIT1 = 16'hf555;
    defparam add_33910_9.INJECT1_0 = "NO";
    defparam add_33910_9.INJECT1_1 = "NO";
    CCU2D add_33910_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48580), .COUT(n48581));
    defparam add_33910_7.INIT0 = 16'hf555;
    defparam add_33910_7.INIT1 = 16'hf555;
    defparam add_33910_7.INJECT1_0 = "NO";
    defparam add_33910_7.INJECT1_1 = "NO";
    PFUMX i38905 (.BLUT(n54895), .ALUT(n54896), .C0(state[1]), .Z(state_2__N_104[2]));
    CCU2D add_33910_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48579), .COUT(n48580));
    defparam add_33910_5.INIT0 = 16'hf555;
    defparam add_33910_5.INIT1 = 16'hf555;
    defparam add_33910_5.INJECT1_0 = "NO";
    defparam add_33910_5.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47803), .COUT(n47804), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47802), .COUT(n47803), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_33910_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48578), .COUT(n48579));
    defparam add_33910_3.INIT0 = 16'hf555;
    defparam add_33910_3.INIT1 = 16'hf555;
    defparam add_33910_3.INJECT1_0 = "NO";
    defparam add_33910_3.INJECT1_1 = "NO";
    CCU2D add_33910_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48578));
    defparam add_33910_1.INIT0 = 16'hF000;
    defparam add_33910_1.INIT1 = 16'ha666;
    defparam add_33910_1.INJECT1_0 = "NO";
    defparam add_33910_1.INJECT1_1 = "NO";
    L6MUX21 i37892 (.D0(n53094), .D1(n53095), .SD(bit_counter[2]), .Z(n53098));
    L6MUX21 i37893 (.D0(n53096), .D1(n53097), .SD(bit_counter[2]), .Z(n53099));
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47801), .COUT(n47802), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47800), .COUT(n47801), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47799), .COUT(n47800), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47798), .COUT(n47799), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47798), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i37711_3_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .D(n13661), .Z(sclk_c_enable_110)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i37711_3_lut_4_lut_4_lut.init = 16'hffc2;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47796), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47795), .COUT(n47796), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47794), .COUT(n47795), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    LUT4 i2459_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n13661), 
         .D(state[0]), .Z(n8556)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2459_4_lut_4_lut_4_lut.init = 16'he8c8;
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47793), .COUT(n47794), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut_then_2_lut (.A(state[2]), .B(n13661), .Z(n55533)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_then_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[7]), 
         .D(state[1]), .Z(n54929)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_then_4_lut.init = 16'hf0f4;
    LUT4 i19509_1_lut_rep_783 (.A(state[2]), .Z(n54786)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i19509_1_lut_rep_783.init = 16'h5555;
    LUT4 i28800_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28800_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_3_lut_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[7]), 
         .D(state[1]), .Z(n54928)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_else_4_lut.init = 16'hf0b0;
    LUT4 mux_2468_i5_4_lut_4_lut_then_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13661), .Z(n54935)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2468_i5_4_lut_4_lut_then_4_lut.init = 16'he2e0;
    LUT4 mux_2468_i5_4_lut_4_lut_else_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13661), .Z(n54934)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2468_i5_4_lut_4_lut_else_4_lut.init = 16'hd0f0;
    LUT4 i1_2_lut_rep_843 (.A(n13626), .B(n11), .Z(n55538)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_843.init = 16'h8888;
    LUT4 i28778_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28778_2_lut.init = 16'hbbbb;
    LUT4 i28777_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_898)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28777_2_lut.init = 16'hbbbb;
    LUT4 mux_2468_i3_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13661), .Z(n54993)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2468_i3_4_lut_then_4_lut.init = 16'hb1f0;
    LUT4 mux_2468_i3_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13626), .Z(n54992)) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2468_i3_4_lut_else_4_lut.init = 16'hb0f4;
    LUT4 i1_2_lut_rep_597_3_lut (.A(state[2]), .B(n13661), .C(state[1]), 
         .Z(n54600)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_597_3_lut.init = 16'h4040;
    LUT4 i38592_3_lut_rep_598_4_lut (.A(state[2]), .B(n13661), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2315)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38592_3_lut_rep_598_4_lut.init = 16'hfffb;
    LUT4 mux_2462_i9_3_lut_4_lut (.A(n13626), .B(n11), .C(n54717), .D(n447[8]), 
         .Z(n8570[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2462_i9_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2462_i10_3_lut_4_lut (.A(n13626), .B(n11), .C(n54717), .D(n447[9]), 
         .Z(n8570[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2462_i10_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2462_i13_3_lut_4_lut (.A(n13626), .B(n11), .C(n54717), .D(n447[12]), 
         .Z(n8570[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2462_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 i30397_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42570)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i30397_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i28709_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15065[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28709_2_lut_3_lut.init = 16'h7070;
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47793), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_714_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54717)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_714_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(n447[0]), 
         .D(state[0]), .Z(n45)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_3_lut_rep_734_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_2133)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_734_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut_adj_133 (.A(state[2]), .B(state[1]), .C(n447[1]), 
         .D(state[0]), .Z(n53)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_133.init = 16'he0f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13661), 
         .Z(sclk_c_enable_106)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_3_lut_4_lut_4_lut_else_2_lut_4_lut (.A(n13626), .B(n11), .C(state[0]), 
         .D(state[2]), .Z(n55532)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_else_2_lut_4_lut.init = 16'h0070;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13626), 
         .D(state[1]), .Z(sclk_c_enable_2100)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_134 (.A(state[0]), .B(state[2]), .C(n13626), 
         .D(state[1]), .Z(n38570)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_134.init = 16'h0002;
    L6MUX21 i38113 (.D0(n53317), .D1(n53318), .SD(bit_counter[2]), .Z(n53319));
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_135 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_135.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_136 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_136.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_137 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_137.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_138 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_138.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_139 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_139.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_140 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_140.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_141 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_141.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_142 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_142.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_143 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_143.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_144 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_144.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_145 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_145.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_146 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_146.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_147 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_147.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_148 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_148.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_149 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_149.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_150 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_150.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_151 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_151.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_152 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_152.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_153 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_153.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_154 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_154.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_155 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_155.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_156 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_156.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_157 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_157.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_158 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_158.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_159 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_159.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_160 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_160.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_161 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_161.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_162 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_162.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_163 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_163.init = 16'h2020;
    LUT4 mux_2452_i2_4_lut_4_lut (.A(n54591), .B(n54717), .C(n8556), .D(n13626), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2452_i2_4_lut_4_lut.init = 16'h5053;
    FD1P3AX delay_counter_i0_i1 (.D(n8746[1]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n8746[3]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n8746[7]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n8746[8]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n8746[9]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n8746[12]), .SP(sclk_c_enable_2315), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3IX pixel_i0 (.D(\Q[11] [0]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i38396_2_lut_rep_829 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_2164)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38396_2_lut_rep_829.init = 16'h9999;
    LUT4 i23542_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35783)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23542_2_lut_2_lut.init = 16'h8888;
    LUT4 i23413_4_lut (.A(sclk_c_enable_2315), .B(n54600), .C(n8745), 
         .D(n54717), .Z(n35605)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23413_4_lut.init = 16'ha8aa;
    PFUMX i37888 (.BLUT(n53086), .ALUT(n53087), .C0(bit_counter[1]), .Z(n53094));
    PFUMX i37889 (.BLUT(n53088), .ALUT(n53089), .C0(bit_counter[1]), .Z(n53095));
    PFUMX i37890 (.BLUT(n53090), .ALUT(n53091), .C0(bit_counter[1]), .Z(n53096));
    PFUMX i37891 (.BLUT(n53092), .ALUT(n53093), .C0(bit_counter[1]), .Z(n53097));
    LUT4 i28931_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i28931_2_lut_3_lut.init = 16'h1010;
    LUT4 i29958_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[8]), .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29958_2_lut_3_lut.init = 16'h1010;
    LUT4 i29962_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[7]), .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29962_2_lut_3_lut.init = 16'h1010;
    LUT4 i29967_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[6]), .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29967_2_lut_3_lut.init = 16'h1010;
    LUT4 i29979_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[5]), .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29979_2_lut_3_lut.init = 16'h1010;
    LUT4 i29986_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[4]), .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29986_2_lut_3_lut.init = 16'h1010;
    LUT4 i29994_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[3]), .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29994_2_lut_3_lut.init = 16'h1010;
    LUT4 i29997_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[2]), .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29997_2_lut_3_lut.init = 16'h1010;
    LUT4 i29998_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[1]), .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29998_2_lut_3_lut.init = 16'h1010;
    LUT4 i38110_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38110_3_lut.init = 16'hcaca;
    LUT4 i38109_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38109_3_lut.init = 16'hcaca;
    LUT4 i38108_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38108_3_lut.init = 16'hcaca;
    LUT4 i38107_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38107_3_lut.init = 16'hcaca;
    LUT4 mux_2478_i1_4_lut (.A(n45), .B(n15065[0]), .C(n8745), .D(n52739), 
         .Z(n8746[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i1_4_lut.init = 16'hcfca;
    LUT4 i2490_3_lut (.A(state[2]), .B(state[1]), .C(n13661), .Z(n8745)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2490_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[6]), .C(n14), .D(cur_pixel[1]), 
         .Z(n11)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[0]), .B(cur_pixel[2]), .C(cur_pixel[8]), 
         .D(cur_pixel[5]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i37887_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37887_3_lut.init = 16'hcaca;
    LUT4 i5_3_lut (.A(cur_pixel[3]), .B(cur_pixel[7]), .C(cur_pixel[4]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i37886_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37886_3_lut.init = 16'hcaca;
    LUT4 i37885_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37885_3_lut.init = 16'hcaca;
    LUT4 i37884_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37884_3_lut.init = 16'hcaca;
    LUT4 i37883_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37883_3_lut.init = 16'hcaca;
    LUT4 i37882_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37882_3_lut.init = 16'hcaca;
    LUT4 i37881_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37881_3_lut.init = 16'hcaca;
    LUT4 i37880_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37880_3_lut.init = 16'hcaca;
    L6MUX21 i37894 (.D0(n53098), .D1(n53099), .SD(bit_counter[3]), .Z(n53100));
    PFUMX i38111 (.BLUT(n53313), .ALUT(n53314), .C0(bit_counter[1]), .Z(n53317));
    PFUMX i38112 (.BLUT(n53315), .ALUT(n53316), .C0(bit_counter[1]), .Z(n53318));
    CCU2D add_3124_33 (.A0(bit_counter[31]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48226), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_33.INIT0 = 16'h5999;
    defparam add_3124_33.INIT1 = 16'h0000;
    defparam add_3124_33.INJECT1_0 = "NO";
    defparam add_3124_33.INJECT1_1 = "NO";
    CCU2D add_33913_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48497), 
          .S0(n13626));
    defparam add_33913_cout.INIT0 = 16'h0000;
    defparam add_33913_cout.INIT1 = 16'h0000;
    defparam add_33913_cout.INJECT1_0 = "NO";
    defparam add_33913_cout.INJECT1_1 = "NO";
    CCU2D add_3124_31 (.A0(bit_counter[29]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48225), .COUT(n48226), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_31.INIT0 = 16'h5999;
    defparam add_3124_31.INIT1 = 16'h5999;
    defparam add_3124_31.INJECT1_0 = "NO";
    defparam add_3124_31.INJECT1_1 = "NO";
    CCU2D add_33913_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48496), .COUT(n48497));
    defparam add_33913_31.INIT0 = 16'hf555;
    defparam add_33913_31.INIT1 = 16'h5555;
    defparam add_33913_31.INJECT1_0 = "NO";
    defparam add_33913_31.INJECT1_1 = "NO";
    CCU2D add_3124_29 (.A0(bit_counter[27]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48224), .COUT(n48225), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_29.INIT0 = 16'h5999;
    defparam add_3124_29.INIT1 = 16'h5999;
    defparam add_3124_29.INJECT1_0 = "NO";
    defparam add_3124_29.INJECT1_1 = "NO";
    CCU2D add_33913_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48495), .COUT(n48496));
    defparam add_33913_29.INIT0 = 16'hf555;
    defparam add_33913_29.INIT1 = 16'hf555;
    defparam add_33913_29.INJECT1_0 = "NO";
    defparam add_33913_29.INJECT1_1 = "NO";
    CCU2D add_3124_27 (.A0(bit_counter[25]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48223), .COUT(n48224), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_27.INIT0 = 16'h5999;
    defparam add_3124_27.INIT1 = 16'h5999;
    defparam add_3124_27.INJECT1_0 = "NO";
    defparam add_3124_27.INJECT1_1 = "NO";
    CCU2D add_33913_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48494), .COUT(n48495));
    defparam add_33913_27.INIT0 = 16'hf555;
    defparam add_33913_27.INIT1 = 16'hf555;
    defparam add_33913_27.INJECT1_0 = "NO";
    defparam add_33913_27.INJECT1_1 = "NO";
    CCU2D add_3124_25 (.A0(bit_counter[23]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48222), .COUT(n48223), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_25.INIT0 = 16'h5999;
    defparam add_3124_25.INIT1 = 16'h5999;
    defparam add_3124_25.INJECT1_0 = "NO";
    defparam add_3124_25.INJECT1_1 = "NO";
    CCU2D add_33913_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48493), .COUT(n48494));
    defparam add_33913_25.INIT0 = 16'hf555;
    defparam add_33913_25.INIT1 = 16'hf555;
    defparam add_33913_25.INJECT1_0 = "NO";
    defparam add_33913_25.INJECT1_1 = "NO";
    CCU2D add_33913_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48492), .COUT(n48493));
    defparam add_33913_23.INIT0 = 16'hf555;
    defparam add_33913_23.INIT1 = 16'hf555;
    defparam add_33913_23.INJECT1_0 = "NO";
    defparam add_33913_23.INJECT1_1 = "NO";
    CCU2D add_3124_23 (.A0(bit_counter[21]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48221), .COUT(n48222), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_23.INIT0 = 16'h5999;
    defparam add_3124_23.INIT1 = 16'h5999;
    defparam add_3124_23.INJECT1_0 = "NO";
    defparam add_3124_23.INJECT1_1 = "NO";
    CCU2D add_3124_21 (.A0(bit_counter[19]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48220), .COUT(n48221), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_21.INIT0 = 16'h5999;
    defparam add_3124_21.INIT1 = 16'h5999;
    defparam add_3124_21.INJECT1_0 = "NO";
    defparam add_3124_21.INJECT1_1 = "NO";
    CCU2D add_3124_19 (.A0(bit_counter[17]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48219), .COUT(n48220), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_19.INIT0 = 16'h5999;
    defparam add_3124_19.INIT1 = 16'h5999;
    defparam add_3124_19.INJECT1_0 = "NO";
    defparam add_3124_19.INJECT1_1 = "NO";
    CCU2D add_3124_17 (.A0(bit_counter[15]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48218), .COUT(n48219), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_17.INIT0 = 16'h5999;
    defparam add_3124_17.INIT1 = 16'h5999;
    defparam add_3124_17.INJECT1_0 = "NO";
    defparam add_3124_17.INJECT1_1 = "NO";
    CCU2D add_33913_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48491), .COUT(n48492));
    defparam add_33913_21.INIT0 = 16'hf555;
    defparam add_33913_21.INIT1 = 16'hf555;
    defparam add_33913_21.INJECT1_0 = "NO";
    defparam add_33913_21.INJECT1_1 = "NO";
    CCU2D add_33913_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48490), .COUT(n48491));
    defparam add_33913_19.INIT0 = 16'hf555;
    defparam add_33913_19.INIT1 = 16'hf555;
    defparam add_33913_19.INJECT1_0 = "NO";
    defparam add_33913_19.INJECT1_1 = "NO";
    CCU2D add_33913_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48489), .COUT(n48490));
    defparam add_33913_17.INIT0 = 16'hf555;
    defparam add_33913_17.INIT1 = 16'hf555;
    defparam add_33913_17.INJECT1_0 = "NO";
    defparam add_33913_17.INJECT1_1 = "NO";
    CCU2D add_33913_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48488), .COUT(n48489));
    defparam add_33913_15.INIT0 = 16'hf555;
    defparam add_33913_15.INIT1 = 16'hf555;
    defparam add_33913_15.INJECT1_0 = "NO";
    defparam add_33913_15.INJECT1_1 = "NO";
    CCU2D add_33913_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48487), .COUT(n48488));
    defparam add_33913_13.INIT0 = 16'hf555;
    defparam add_33913_13.INIT1 = 16'hf555;
    defparam add_33913_13.INJECT1_0 = "NO";
    defparam add_33913_13.INJECT1_1 = "NO";
    CCU2D add_3124_15 (.A0(bit_counter[13]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48217), .COUT(n48218), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_15.INIT0 = 16'h5999;
    defparam add_3124_15.INIT1 = 16'h5999;
    defparam add_3124_15.INJECT1_0 = "NO";
    defparam add_3124_15.INJECT1_1 = "NO";
    CCU2D add_3124_13 (.A0(bit_counter[11]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48216), .COUT(n48217), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_13.INIT0 = 16'h5999;
    defparam add_3124_13.INIT1 = 16'h5999;
    defparam add_3124_13.INJECT1_0 = "NO";
    defparam add_3124_13.INJECT1_1 = "NO";
    CCU2D add_3124_11 (.A0(bit_counter[9]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48215), .COUT(n48216), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_11.INIT0 = 16'h5999;
    defparam add_3124_11.INIT1 = 16'h5999;
    defparam add_3124_11.INJECT1_0 = "NO";
    defparam add_3124_11.INJECT1_1 = "NO";
    CCU2D add_3124_9 (.A0(bit_counter[7]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48214), .COUT(n48215), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_9.INIT0 = 16'h5999;
    defparam add_3124_9.INIT1 = 16'h5999;
    defparam add_3124_9.INJECT1_0 = "NO";
    defparam add_3124_9.INJECT1_1 = "NO";
    CCU2D add_3124_7 (.A0(bit_counter[5]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48213), .COUT(n48214), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_7.INIT0 = 16'h5999;
    defparam add_3124_7.INIT1 = 16'h5999;
    defparam add_3124_7.INJECT1_0 = "NO";
    defparam add_3124_7.INJECT1_1 = "NO";
    CCU2D add_3124_5 (.A0(bit_counter[3]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48212), .COUT(n48213), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_5.INIT0 = 16'h5999;
    defparam add_3124_5.INIT1 = 16'h5999;
    defparam add_3124_5.INJECT1_0 = "NO";
    defparam add_3124_5.INJECT1_1 = "NO";
    CCU2D add_3124_3 (.A0(bit_counter[1]), .B0(n13626), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13626), .C1(GND_net), 
          .D1(GND_net), .CIN(n48211), .COUT(n48212), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_3.INIT0 = 16'h5999;
    defparam add_3124_3.INIT1 = 16'h5999;
    defparam add_3124_3.INJECT1_0 = "NO";
    defparam add_3124_3.INJECT1_1 = "NO";
    CCU2D add_33913_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48486), .COUT(n48487));
    defparam add_33913_11.INIT0 = 16'hf555;
    defparam add_33913_11.INIT1 = 16'hf555;
    defparam add_33913_11.INJECT1_0 = "NO";
    defparam add_33913_11.INJECT1_1 = "NO";
    CCU2D add_3124_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13626), .C1(GND_net), .D1(GND_net), 
          .COUT(n48211), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3124_1.INIT0 = 16'hF000;
    defparam add_3124_1.INIT1 = 16'h5999;
    defparam add_3124_1.INJECT1_0 = "NO";
    defparam add_3124_1.INJECT1_1 = "NO";
    CCU2D add_33913_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48485), .COUT(n48486));
    defparam add_33913_9.INIT0 = 16'hf555;
    defparam add_33913_9.INIT1 = 16'hf555;
    defparam add_33913_9.INJECT1_0 = "NO";
    defparam add_33913_9.INJECT1_1 = "NO";
    CCU2D add_33913_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48484), .COUT(n48485));
    defparam add_33913_7.INIT0 = 16'hf555;
    defparam add_33913_7.INIT1 = 16'hf555;
    defparam add_33913_7.INJECT1_0 = "NO";
    defparam add_33913_7.INJECT1_1 = "NO";
    CCU2D add_33913_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48483), .COUT(n48484));
    defparam add_33913_5.INIT0 = 16'hf555;
    defparam add_33913_5.INIT1 = 16'hf555;
    defparam add_33913_5.INJECT1_0 = "NO";
    defparam add_33913_5.INJECT1_1 = "NO";
    CCU2D add_33913_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48482), .COUT(n48483));
    defparam add_33913_3.INIT0 = 16'hf555;
    defparam add_33913_3.INIT1 = 16'hf555;
    defparam add_33913_3.INJECT1_0 = "NO";
    defparam add_33913_3.INJECT1_1 = "NO";
    CCU2D add_33913_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48482));
    defparam add_33913_1.INIT0 = 16'hF000;
    defparam add_33913_1.INIT1 = 16'ha666;
    defparam add_33913_1.INJECT1_0 = "NO";
    defparam add_33913_1.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53100), .B(n53319), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 mux_2452_i1_4_lut (.A(n54717), .B(n54591), .C(n8556), .D(n55538), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2452_i1_4_lut.init = 16'h3f3a;
    FD1P3IX pixel_i23 (.D(\Q[11] [23]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[11] [22]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[11] [21]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[11] [20]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[11] [19]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[11] [18]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[11] [17]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[11] [16]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[11] [15]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[11] [14]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[11] [13]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[11] [12]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[11] [11]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[11] [10]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[11] [9]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[11] [8]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[11] [7]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[11] [6]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[11] [5]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[11] [4]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[11] [3]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[11] [2]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[11] [1]), .SP(sclk_c_enable_2133), .CD(n35783), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2100), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2133), 
            .CD(n35783), .CK(sclk_c), .Q(\RdAddress[11] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_2164), .CD(n35783), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_898), .SP(sclk_c_enable_2164), .CD(n35783), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_2164), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2315), 
            .CD(n35605), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2315), .CD(n35605), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2315), .CD(n35605), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54936), .SP(sclk_c_enable_2315), .CD(n8745), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54994), .SP(sclk_c_enable_2315), .CD(n8745), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=256, LSE_RLINE=256 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 mux_2452_i3_4_lut_then_3_lut (.A(state[0]), .B(n13661), .C(state[2]), 
         .Z(n54896)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2452_i3_4_lut_then_3_lut.init = 16'h0808;
    LUT4 mux_2478_i2_4_lut (.A(n53), .B(n15065[0]), .C(n8745), .D(n52739), 
         .Z(n8746[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2478_i4_4_lut (.A(n38570), .B(n42570), .C(n8745), .D(n4), 
         .Z(n8746[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n11), .B(n54600), .C(n447[3]), .D(n54717), .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 mux_2478_i8_4_lut (.A(n54930), .B(n42570), .C(n8745), .D(n54600), 
         .Z(n8746[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i8_4_lut.init = 16'h303a;
    LUT4 mux_2478_i9_4_lut (.A(n8570[8]), .B(n42570), .C(n8745), .D(n54600), 
         .Z(n8746[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i9_4_lut.init = 16'h303a;
    LUT4 mux_2478_i10_4_lut (.A(n8570[9]), .B(n42570), .C(n8745), .D(n54600), 
         .Z(n8746[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i10_4_lut.init = 16'h303a;
    LUT4 mux_2478_i13_4_lut (.A(n8570[12]), .B(n42570), .C(n8745), .D(n54600), 
         .Z(n8746[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2478_i13_4_lut.init = 16'h303a;
    LUT4 mux_2452_i3_4_lut_else_3_lut (.A(state[0]), .B(state[2]), .C(n11), 
         .D(n13626), .Z(n54895)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2452_i3_4_lut_else_3_lut.init = 16'h2000;
    PFUMX i38969 (.BLUT(n54992), .ALUT(n54993), .C0(state[1]), .Z(n54994));
    PFUMX i38931 (.BLUT(n54934), .ALUT(n54935), .C0(state[0]), .Z(n54936));
    PFUMX i39241 (.BLUT(n55532), .ALUT(n55533), .C0(state[1]), .Z(n52739));
    PFUMX i38927 (.BLUT(n54928), .ALUT(n54929), .C0(n55538), .Z(n54930));
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47813), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47812), .COUT(n47813), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47811), .COUT(n47812), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_33910_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48593), 
          .S0(n13661));
    defparam add_33910_cout.INIT0 = 16'h0000;
    defparam add_33910_cout.INIT1 = 16'h0000;
    defparam add_33910_cout.INJECT1_0 = "NO";
    defparam add_33910_cout.INJECT1_1 = "NO";
    CCU2D add_33910_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48592), .COUT(n48593));
    defparam add_33910_31.INIT0 = 16'hf555;
    defparam add_33910_31.INIT1 = 16'h5555;
    defparam add_33910_31.INJECT1_0 = "NO";
    defparam add_33910_31.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47810), .COUT(n47811), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47809), .COUT(n47810), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47808), .COUT(n47809), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_33910_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48591), .COUT(n48592));
    defparam add_33910_29.INIT0 = 16'hf555;
    defparam add_33910_29.INIT1 = 16'hf555;
    defparam add_33910_29.INJECT1_0 = "NO";
    defparam add_33910_29.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47807), .COUT(n47808), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_33910_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48590), .COUT(n48591));
    defparam add_33910_27.INIT0 = 16'hf555;
    defparam add_33910_27.INIT1 = 16'hf555;
    defparam add_33910_27.INJECT1_0 = "NO";
    defparam add_33910_27.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47806), .COUT(n47807), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47805), .COUT(n47806), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_33910_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48589), .COUT(n48590));
    defparam add_33910_25.INIT0 = 16'hf555;
    defparam add_33910_25.INIT1 = 16'hf555;
    defparam add_33910_25.INJECT1_0 = "NO";
    defparam add_33910_25.INJECT1_1 = "NO";
    CCU2D add_33910_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48588), .COUT(n48589));
    defparam add_33910_23.INIT0 = 16'hf555;
    defparam add_33910_23.INIT1 = 16'hf555;
    defparam add_33910_23.INJECT1_0 = "NO";
    defparam add_33910_23.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U38 
//

module \WS2812(48000000,"111111111")_U38  (sclk_c, \port_status[10] , ws2813_out_c_10, 
            GND_net, \Q[10] , \RdAddress[10] );
    input sclk_c;
    output \port_status[10] ;
    output ws2813_out_c_10;
    input GND_net;
    input [23:0]\Q[10] ;
    output [8:0]\RdAddress[10] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire n42702, n13556, n54637;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_2410;
    wire [31:0]n8479;
    
    wire sclk_c_enable_94, n54791, sclk_c_enable_95, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_98;
    wire [2:0]state_2__N_104;
    
    wire n53079, n53080;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53083, n53081, n53082, n53084;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire n15, n54594, n13591, sclk_c_enable_2195, n54902, n54901, 
        n54648, n54743, serial_N_437;
    wire [31:0]n447;
    
    wire n54978, n54977, n54721;
    wire [31:0]n8303;
    
    wire n80, n14, n53310, n53311, n53312, n47792, n47791;
    wire [6:0]n15057;
    
    wire n42564, n54809, n71, sclk_c_enable_2228, n74, n35688;
    wire [31:0]bit_counter_31__N_204;
    
    wire n1, n1_adj_897;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    wire [8:0]cur_pixel_8__N_107;
    
    wire sclk_c_enable_2259;
    wire [31:0]bit_counter_31__N_172;
    
    wire n35659, n47790, n47789, n47788, n47787, n47786, n47785, 
        n47784, n47783, n53071, n53072, n47782, n53073, n53074, 
        n53075, n53076, n53077, n53078, n47781, n47780, n47779, 
        n47778, n47777;
    wire [8:0]n118;
    
    wire n54620, n52742, n53309, n53308, n53307, n53306, n8478, 
        n54579, n35510, n47775, n35506, n48258, n48257, n48256, 
        n47774;
    wire [2:0]n8806;
    wire [31:0]n8405;
    
    wire n47773, n48255, n48254, n48253, n48252, n48251, n47772, 
        n48250, n48249, n48248, n53085, n48247, n48246, n48245, 
        n48244, n48243, n38671, n48481, n48480, n48479, n48478, 
        n48477, n48476, n48475, n48474, n48473, n48472, n48471, 
        n48470, n48469, n48468, n48467, n48466, n48465, n48464, 
        n48463, n48462, n48461, n8813, n48460, n48459, n48458, 
        n48457, n48456, n48455, n48454, n48453, n48452, n48451, 
        n48450, n54979, n4;
    
    LUT4 i37687_2_lut_rep_634 (.A(n42702), .B(n13556), .Z(n54637)) /* synthesis lut_function=(A (B)) */ ;
    defparam i37687_2_lut_rep_634.init = 16'h8888;
    FD1P3AX delay_counter_i0_i0 (.D(n8479[0]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54791), .SP(sclk_c_enable_94), .CK(sclk_c), 
            .Q(\port_status[10] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_95), .CK(sclk_c), 
            .Q(ws2813_out_c_10)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_98), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_98), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_98), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    L6MUX21 i37877 (.D0(n53079), .D1(n53080), .SD(bit_counter[2]), .Z(n53083));
    L6MUX21 i37878 (.D0(n53081), .D1(n53082), .SD(bit_counter[2]), .Z(n53084));
    LUT4 i6_4_lut (.A(cur_pixel[2]), .B(cur_pixel[7]), .C(cur_pixel[5]), 
         .D(cur_pixel[4]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_591_3_lut (.A(n42702), .B(n13556), .C(state[1]), 
         .Z(n54594)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_591_3_lut.init = 16'h0808;
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13591), .Z(sclk_c_enable_98)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n13556), 
         .D(state[0]), .Z(sclk_c_enable_2195)) /* synthesis lut_function=(A (B)+!A !(B+!(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h9888;
    LUT4 i38477_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n13591), 
         .Z(n54902)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38477_4_lut_then_3_lut.init = 16'h1010;
    LUT4 i38477_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n13556), 
         .Z(n54901)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38477_4_lut_else_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_645 (.A(state[1]), .B(n13591), .Z(n54648)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_645.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[1]), .B(n13591), .C(n54743), .D(n54637), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd080;
    LUT4 i21989_1_lut_rep_788 (.A(state[2]), .Z(n54791)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i21989_1_lut_rep_788.init = 16'h5555;
    LUT4 i28805_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28805_3_lut_3_lut.init = 16'h5151;
    LUT4 mux_2411_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13591), .Z(n54978)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2411_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_2411_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13556), .Z(n54977)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2411_i3_4_lut_else_4_lut.init = 16'hd0f2;
    LUT4 i1_3_lut_4_lut (.A(n54594), .B(n54743), .C(n447[7]), .D(n54721), 
         .Z(n8303[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_86 (.A(n54594), .B(n54743), .C(n447[8]), .D(n54721), 
         .Z(n8303[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_86.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_87 (.A(n54594), .B(n54743), .C(n447[9]), .D(n54721), 
         .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_87.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_88 (.A(n54594), .B(n54743), .C(n447[12]), 
         .D(n54721), .Z(n8303[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_88.init = 16'hf888;
    LUT4 i5_3_lut (.A(cur_pixel[8]), .B(cur_pixel[0]), .C(cur_pixel[1]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i5_3_lut.init = 16'h8080;
    L6MUX21 i38106 (.D0(n53310), .D1(n53311), .SD(bit_counter[2]), .Z(n53312));
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47792), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47791), .COUT(n47792), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n15057[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i30392_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42564)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i30392_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_806 (.A(state[1]), .B(state[2]), .Z(n54809)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_806.init = 16'heeee;
    LUT4 i1_2_lut_rep_718_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54721)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_718_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_3_lut_rep_731_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(sclk_c_enable_2228)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_731_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut_adj_89 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_89.init = 16'he0f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(n13591), 
         .Z(sclk_c_enable_95)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i23539_2_lut_4_lut_4_lut_2_lut (.A(state[1]), .B(state[2]), .Z(n35688)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i23539_2_lut_4_lut_4_lut_2_lut.init = 16'h8888;
    FD1P3AX delay_counter_i0_i1 (.D(n8479[1]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n8479[3]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n8479[7]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n8479[8]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n8479[9]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n8479[12]), .SP(sclk_c_enable_2410), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    LUT4 i28776_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28776_2_lut.init = 16'hbbbb;
    LUT4 i28775_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_897)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28775_2_lut.init = 16'hbbbb;
    FD1P3IX pixel_i0 (.D(\Q[10] [0]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i38422_2_lut_rep_827 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_2259)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38422_2_lut_rep_827.init = 16'h9999;
    LUT4 i23447_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35659)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23447_2_lut_2_lut.init = 16'h8888;
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47790), .COUT(n47791), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47789), .COUT(n47790), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47788), .COUT(n47789), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47787), .COUT(n47788), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47786), .COUT(n47787), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47785), .COUT(n47786), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47784), .COUT(n47785), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47783), .COUT(n47784), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    PFUMX i37873 (.BLUT(n53071), .ALUT(n53072), .C0(bit_counter[1]), .Z(n53079));
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47782), .COUT(n47783), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    PFUMX i37874 (.BLUT(n53073), .ALUT(n53074), .C0(bit_counter[1]), .Z(n53080));
    PFUMX i37875 (.BLUT(n53075), .ALUT(n53076), .C0(bit_counter[1]), .Z(n53081));
    PFUMX i37876 (.BLUT(n53077), .ALUT(n53078), .C0(bit_counter[1]), .Z(n53082));
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47781), .COUT(n47782), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47780), .COUT(n47781), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47779), .COUT(n47780), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47778), .COUT(n47779), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47777), .COUT(n47778), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47777), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_90 (.A(state[2]), .B(n42702), .C(n118[0]), 
         .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_90.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_91 (.A(state[2]), .B(n42702), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_91.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_92 (.A(state[2]), .B(n42702), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_92.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_93 (.A(state[2]), .B(n42702), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_93.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_94 (.A(state[2]), .B(n42702), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_94.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_95 (.A(state[2]), .B(n42702), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_95.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_96 (.A(state[2]), .B(n42702), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_96.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_97 (.A(state[2]), .B(n42702), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_97.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_98 (.A(state[2]), .B(n42702), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_98.init = 16'h1010;
    LUT4 i1_3_lut_4_lut_4_lut_adj_99 (.A(n54743), .B(state[1]), .C(n54637), 
         .D(n54620), .Z(n52742)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_99.init = 16'hce02;
    LUT4 i38103_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38103_3_lut.init = 16'hcaca;
    LUT4 i38102_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38102_3_lut.init = 16'hcaca;
    LUT4 i38101_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38101_3_lut.init = 16'hcaca;
    LUT4 i38100_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38100_3_lut.init = 16'hcaca;
    LUT4 i23318_4_lut (.A(sclk_c_enable_2410), .B(n54721), .C(n8478), 
         .D(n54579), .Z(n35510)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23318_4_lut.init = 16'haaa2;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47775), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[6]), .C(n14), .D(cur_pixel[3]), 
         .Z(n42702)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(68[10:33])
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i23294_2_lut_4_lut (.A(n54620), .B(state[0]), .C(state[1]), .D(n8478), 
         .Z(n35506)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23294_2_lut_4_lut.init = 16'hfd00;
    CCU2D add_3122_33 (.A0(bit_counter[31]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48258), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_33.INIT0 = 16'h5999;
    defparam add_3122_33.INIT1 = 16'h0000;
    defparam add_3122_33.INJECT1_0 = "NO";
    defparam add_3122_33.INJECT1_1 = "NO";
    CCU2D add_3122_31 (.A0(bit_counter[29]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48257), .COUT(n48258), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_31.INIT0 = 16'h5999;
    defparam add_3122_31.INIT1 = 16'h5999;
    defparam add_3122_31.INJECT1_0 = "NO";
    defparam add_3122_31.INJECT1_1 = "NO";
    CCU2D add_3122_29 (.A0(bit_counter[27]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48256), .COUT(n48257), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_29.INIT0 = 16'h5999;
    defparam add_3122_29.INIT1 = 16'h5999;
    defparam add_3122_29.INJECT1_0 = "NO";
    defparam add_3122_29.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47774), .COUT(n47775), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_100 (.A(state[0]), .B(n54809), .C(n13556), 
         .D(n42702), .Z(n8806[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_100.init = 16'hfddd;
    LUT4 mux_2411_i5_4_lut_4_lut (.A(state[0]), .B(n54809), .C(n447[4]), 
         .D(n54579), .Z(n8405[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2411_i5_4_lut_4_lut.init = 16'haad0;
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47773), .COUT(n47774), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_3122_27 (.A0(bit_counter[25]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48255), .COUT(n48256), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_27.INIT0 = 16'h5999;
    defparam add_3122_27.INIT1 = 16'h5999;
    defparam add_3122_27.INJECT1_0 = "NO";
    defparam add_3122_27.INJECT1_1 = "NO";
    CCU2D add_3122_25 (.A0(bit_counter[23]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48254), .COUT(n48255), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_25.INIT0 = 16'h5999;
    defparam add_3122_25.INIT1 = 16'h5999;
    defparam add_3122_25.INJECT1_0 = "NO";
    defparam add_3122_25.INJECT1_1 = "NO";
    CCU2D add_3122_23 (.A0(bit_counter[21]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48253), .COUT(n48254), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_23.INIT0 = 16'h5999;
    defparam add_3122_23.INIT1 = 16'h5999;
    defparam add_3122_23.INJECT1_0 = "NO";
    defparam add_3122_23.INJECT1_1 = "NO";
    CCU2D add_3122_21 (.A0(bit_counter[19]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48252), .COUT(n48253), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_21.INIT0 = 16'h5999;
    defparam add_3122_21.INIT1 = 16'h5999;
    defparam add_3122_21.INJECT1_0 = "NO";
    defparam add_3122_21.INJECT1_1 = "NO";
    CCU2D add_3122_19 (.A0(bit_counter[17]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48251), .COUT(n48252), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_19.INIT0 = 16'h5999;
    defparam add_3122_19.INIT1 = 16'h5999;
    defparam add_3122_19.INJECT1_0 = "NO";
    defparam add_3122_19.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47772), .COUT(n47773), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_3122_17 (.A0(bit_counter[15]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48250), .COUT(n48251), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_17.INIT0 = 16'h5999;
    defparam add_3122_17.INIT1 = 16'h5999;
    defparam add_3122_17.INJECT1_0 = "NO";
    defparam add_3122_17.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47772), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    CCU2D add_3122_15 (.A0(bit_counter[13]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48249), .COUT(n48250), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_15.INIT0 = 16'h5999;
    defparam add_3122_15.INIT1 = 16'h5999;
    defparam add_3122_15.INJECT1_0 = "NO";
    defparam add_3122_15.INJECT1_1 = "NO";
    CCU2D add_3122_13 (.A0(bit_counter[11]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48248), .COUT(n48249), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_13.INIT0 = 16'h5999;
    defparam add_3122_13.INIT1 = 16'h5999;
    defparam add_3122_13.INJECT1_0 = "NO";
    defparam add_3122_13.INJECT1_1 = "NO";
    L6MUX21 i37879 (.D0(n53083), .D1(n53084), .SD(bit_counter[3]), .Z(n53085));
    CCU2D add_3122_11 (.A0(bit_counter[9]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48247), .COUT(n48248), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_11.INIT0 = 16'h5999;
    defparam add_3122_11.INIT1 = 16'h5999;
    defparam add_3122_11.INJECT1_0 = "NO";
    defparam add_3122_11.INJECT1_1 = "NO";
    CCU2D add_3122_9 (.A0(bit_counter[7]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48246), .COUT(n48247), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_9.INIT0 = 16'h5999;
    defparam add_3122_9.INIT1 = 16'h5999;
    defparam add_3122_9.INJECT1_0 = "NO";
    defparam add_3122_9.INJECT1_1 = "NO";
    CCU2D add_3122_7 (.A0(bit_counter[5]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48245), .COUT(n48246), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_7.INIT0 = 16'h5999;
    defparam add_3122_7.INIT1 = 16'h5999;
    defparam add_3122_7.INJECT1_0 = "NO";
    defparam add_3122_7.INJECT1_1 = "NO";
    LUT4 i37872_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37872_3_lut.init = 16'hcaca;
    LUT4 i37871_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37871_3_lut.init = 16'hcaca;
    LUT4 i37870_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37870_3_lut.init = 16'hcaca;
    LUT4 i37869_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37869_3_lut.init = 16'hcaca;
    LUT4 i37868_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37868_3_lut.init = 16'hcaca;
    LUT4 i37867_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37867_3_lut.init = 16'hcaca;
    LUT4 i37866_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37866_3_lut.init = 16'hcaca;
    LUT4 i37865_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37865_3_lut.init = 16'hcaca;
    CCU2D add_3122_5 (.A0(bit_counter[3]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48244), .COUT(n48245), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_5.INIT0 = 16'h5999;
    defparam add_3122_5.INIT1 = 16'h5999;
    defparam add_3122_5.INJECT1_0 = "NO";
    defparam add_3122_5.INJECT1_1 = "NO";
    CCU2D add_3122_3 (.A0(bit_counter[1]), .B0(n13556), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13556), .C1(GND_net), 
          .D1(GND_net), .CIN(n48243), .COUT(n48244), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_3.INIT0 = 16'h5999;
    defparam add_3122_3.INIT1 = 16'h5999;
    defparam add_3122_3.INJECT1_0 = "NO";
    defparam add_3122_3.INJECT1_1 = "NO";
    CCU2D add_3122_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13556), .C1(GND_net), .D1(GND_net), 
          .COUT(n48243), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3122_1.INIT0 = 16'hF000;
    defparam add_3122_1.INIT1 = 16'h5999;
    defparam add_3122_1.INJECT1_0 = "NO";
    defparam add_3122_1.INJECT1_1 = "NO";
    PFUMX i38104 (.BLUT(n53306), .ALUT(n53307), .C0(bit_counter[1]), .Z(n53310));
    PFUMX i38105 (.BLUT(n53308), .ALUT(n53309), .C0(bit_counter[1]), .Z(n53311));
    LUT4 i1_2_lut_rep_740 (.A(state[2]), .B(state[0]), .Z(n54743)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_740.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_101 (.A(state[2]), .B(state[0]), .C(n13556), 
         .D(state[1]), .Z(n38671)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_101.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_adj_102 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_102.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_103 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_103.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_104 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_104.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_105 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_105.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_106 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_106.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_107 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_107.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_108 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_108.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_109 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_109.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_110 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_110.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_111 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_111.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_112 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_112.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_113 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_113.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_114 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_114.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_115 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_115.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_116 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_116.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_117 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_117.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_118 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_118.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_119 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_119.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_120 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_120.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_121 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_121.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_122 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_122.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_123 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_123.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_124 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_124.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_125 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_125.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_126 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_126.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_127 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_127.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_128 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_128.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_129 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_129.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_130 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_130.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_131 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_131.init = 16'h4040;
    CCU2D add_33914_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48481), 
          .S0(n13591));
    defparam add_33914_cout.INIT0 = 16'h0000;
    defparam add_33914_cout.INIT1 = 16'h0000;
    defparam add_33914_cout.INJECT1_0 = "NO";
    defparam add_33914_cout.INJECT1_1 = "NO";
    CCU2D add_33914_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48480), .COUT(n48481));
    defparam add_33914_31.INIT0 = 16'hf555;
    defparam add_33914_31.INIT1 = 16'h5555;
    defparam add_33914_31.INJECT1_0 = "NO";
    defparam add_33914_31.INJECT1_1 = "NO";
    CCU2D add_33914_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48479), .COUT(n48480));
    defparam add_33914_29.INIT0 = 16'hf555;
    defparam add_33914_29.INIT1 = 16'hf555;
    defparam add_33914_29.INJECT1_0 = "NO";
    defparam add_33914_29.INJECT1_1 = "NO";
    CCU2D add_33914_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48478), .COUT(n48479));
    defparam add_33914_27.INIT0 = 16'hf555;
    defparam add_33914_27.INIT1 = 16'hf555;
    defparam add_33914_27.INJECT1_0 = "NO";
    defparam add_33914_27.INJECT1_1 = "NO";
    CCU2D add_33914_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48477), .COUT(n48478));
    defparam add_33914_25.INIT0 = 16'hf555;
    defparam add_33914_25.INIT1 = 16'hf555;
    defparam add_33914_25.INJECT1_0 = "NO";
    defparam add_33914_25.INJECT1_1 = "NO";
    CCU2D add_33914_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48476), .COUT(n48477));
    defparam add_33914_23.INIT0 = 16'hf555;
    defparam add_33914_23.INIT1 = 16'hf555;
    defparam add_33914_23.INJECT1_0 = "NO";
    defparam add_33914_23.INJECT1_1 = "NO";
    CCU2D add_33914_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48475), .COUT(n48476));
    defparam add_33914_21.INIT0 = 16'hf555;
    defparam add_33914_21.INIT1 = 16'hf555;
    defparam add_33914_21.INJECT1_0 = "NO";
    defparam add_33914_21.INJECT1_1 = "NO";
    CCU2D add_33914_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48474), .COUT(n48475));
    defparam add_33914_19.INIT0 = 16'hf555;
    defparam add_33914_19.INIT1 = 16'hf555;
    defparam add_33914_19.INJECT1_0 = "NO";
    defparam add_33914_19.INJECT1_1 = "NO";
    CCU2D add_33914_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48473), .COUT(n48474));
    defparam add_33914_17.INIT0 = 16'hf555;
    defparam add_33914_17.INIT1 = 16'hf555;
    defparam add_33914_17.INJECT1_0 = "NO";
    defparam add_33914_17.INJECT1_1 = "NO";
    CCU2D add_33914_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48472), .COUT(n48473));
    defparam add_33914_15.INIT0 = 16'hf555;
    defparam add_33914_15.INIT1 = 16'hf555;
    defparam add_33914_15.INJECT1_0 = "NO";
    defparam add_33914_15.INJECT1_1 = "NO";
    CCU2D add_33914_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48471), .COUT(n48472));
    defparam add_33914_13.INIT0 = 16'hf555;
    defparam add_33914_13.INIT1 = 16'hf555;
    defparam add_33914_13.INJECT1_0 = "NO";
    defparam add_33914_13.INJECT1_1 = "NO";
    CCU2D add_33914_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48470), .COUT(n48471));
    defparam add_33914_11.INIT0 = 16'hf555;
    defparam add_33914_11.INIT1 = 16'hf555;
    defparam add_33914_11.INJECT1_0 = "NO";
    defparam add_33914_11.INJECT1_1 = "NO";
    CCU2D add_33914_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48469), .COUT(n48470));
    defparam add_33914_9.INIT0 = 16'hf555;
    defparam add_33914_9.INIT1 = 16'hf555;
    defparam add_33914_9.INJECT1_0 = "NO";
    defparam add_33914_9.INJECT1_1 = "NO";
    CCU2D add_33914_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48468), .COUT(n48469));
    defparam add_33914_7.INIT0 = 16'hf555;
    defparam add_33914_7.INIT1 = 16'hf555;
    defparam add_33914_7.INJECT1_0 = "NO";
    defparam add_33914_7.INJECT1_1 = "NO";
    CCU2D add_33914_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48467), .COUT(n48468));
    defparam add_33914_5.INIT0 = 16'hf555;
    defparam add_33914_5.INIT1 = 16'hf555;
    defparam add_33914_5.INJECT1_0 = "NO";
    defparam add_33914_5.INJECT1_1 = "NO";
    CCU2D add_33914_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48466), .COUT(n48467));
    defparam add_33914_3.INIT0 = 16'hf555;
    defparam add_33914_3.INIT1 = 16'hf555;
    defparam add_33914_3.INJECT1_0 = "NO";
    defparam add_33914_3.INJECT1_1 = "NO";
    CCU2D add_33914_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48466));
    defparam add_33914_1.INIT0 = 16'hF000;
    defparam add_33914_1.INIT1 = 16'ha666;
    defparam add_33914_1.INJECT1_0 = "NO";
    defparam add_33914_1.INJECT1_1 = "NO";
    CCU2D add_33915_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48465), 
          .S0(n13556));
    defparam add_33915_cout.INIT0 = 16'h0000;
    defparam add_33915_cout.INIT1 = 16'h0000;
    defparam add_33915_cout.INJECT1_0 = "NO";
    defparam add_33915_cout.INJECT1_1 = "NO";
    CCU2D add_33915_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48464), .COUT(n48465));
    defparam add_33915_31.INIT0 = 16'hf555;
    defparam add_33915_31.INIT1 = 16'h5555;
    defparam add_33915_31.INJECT1_0 = "NO";
    defparam add_33915_31.INJECT1_1 = "NO";
    CCU2D add_33915_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48463), .COUT(n48464));
    defparam add_33915_29.INIT0 = 16'hf555;
    defparam add_33915_29.INIT1 = 16'hf555;
    defparam add_33915_29.INJECT1_0 = "NO";
    defparam add_33915_29.INJECT1_1 = "NO";
    CCU2D add_33915_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48462), .COUT(n48463));
    defparam add_33915_27.INIT0 = 16'hf555;
    defparam add_33915_27.INIT1 = 16'hf555;
    defparam add_33915_27.INJECT1_0 = "NO";
    defparam add_33915_27.INJECT1_1 = "NO";
    CCU2D add_33915_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48461), .COUT(n48462));
    defparam add_33915_25.INIT0 = 16'hf555;
    defparam add_33915_25.INIT1 = 16'hf555;
    defparam add_33915_25.INJECT1_0 = "NO";
    defparam add_33915_25.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53085), .B(n53312), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i29567_4_lut (.A(n8806[0]), .B(n8813), .C(state[0]), .D(n54648), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29567_4_lut.init = 16'h0322;
    LUT4 i1_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(n13591), 
         .Z(n8813)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut.init = 16'ha8a0;
    CCU2D add_33915_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48460), .COUT(n48461));
    defparam add_33915_23.INIT0 = 16'hf555;
    defparam add_33915_23.INIT1 = 16'hf555;
    defparam add_33915_23.INJECT1_0 = "NO";
    defparam add_33915_23.INJECT1_1 = "NO";
    CCU2D add_33915_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48459), .COUT(n48460));
    defparam add_33915_21.INIT0 = 16'hf555;
    defparam add_33915_21.INIT1 = 16'hf555;
    defparam add_33915_21.INJECT1_0 = "NO";
    defparam add_33915_21.INJECT1_1 = "NO";
    CCU2D add_33915_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48458), .COUT(n48459));
    defparam add_33915_19.INIT0 = 16'hf555;
    defparam add_33915_19.INIT1 = 16'hf555;
    defparam add_33915_19.INJECT1_0 = "NO";
    defparam add_33915_19.INJECT1_1 = "NO";
    CCU2D add_33915_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48457), .COUT(n48458));
    defparam add_33915_17.INIT0 = 16'hf555;
    defparam add_33915_17.INIT1 = 16'hf555;
    defparam add_33915_17.INJECT1_0 = "NO";
    defparam add_33915_17.INJECT1_1 = "NO";
    CCU2D add_33915_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48456), .COUT(n48457));
    defparam add_33915_15.INIT0 = 16'hf555;
    defparam add_33915_15.INIT1 = 16'hf555;
    defparam add_33915_15.INJECT1_0 = "NO";
    defparam add_33915_15.INJECT1_1 = "NO";
    CCU2D add_33915_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48455), .COUT(n48456));
    defparam add_33915_13.INIT0 = 16'hf555;
    defparam add_33915_13.INIT1 = 16'hf555;
    defparam add_33915_13.INJECT1_0 = "NO";
    defparam add_33915_13.INJECT1_1 = "NO";
    CCU2D add_33915_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48454), .COUT(n48455));
    defparam add_33915_11.INIT0 = 16'hf555;
    defparam add_33915_11.INIT1 = 16'hf555;
    defparam add_33915_11.INJECT1_0 = "NO";
    defparam add_33915_11.INJECT1_1 = "NO";
    CCU2D add_33915_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48453), .COUT(n48454));
    defparam add_33915_9.INIT0 = 16'hf555;
    defparam add_33915_9.INIT1 = 16'hf555;
    defparam add_33915_9.INJECT1_0 = "NO";
    defparam add_33915_9.INJECT1_1 = "NO";
    CCU2D add_33915_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48452), .COUT(n48453));
    defparam add_33915_7.INIT0 = 16'hf555;
    defparam add_33915_7.INIT1 = 16'hf555;
    defparam add_33915_7.INJECT1_0 = "NO";
    defparam add_33915_7.INJECT1_1 = "NO";
    CCU2D add_33915_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48451), .COUT(n48452));
    defparam add_33915_5.INIT0 = 16'hf555;
    defparam add_33915_5.INIT1 = 16'hf555;
    defparam add_33915_5.INJECT1_0 = "NO";
    defparam add_33915_5.INJECT1_1 = "NO";
    CCU2D add_33915_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48450), .COUT(n48451));
    defparam add_33915_3.INIT0 = 16'hf555;
    defparam add_33915_3.INIT1 = 16'hf555;
    defparam add_33915_3.INJECT1_0 = "NO";
    defparam add_33915_3.INJECT1_1 = "NO";
    CCU2D add_33915_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48450));
    defparam add_33915_1.INIT0 = 16'hF000;
    defparam add_33915_1.INIT1 = 16'ha666;
    defparam add_33915_1.INJECT1_0 = "NO";
    defparam add_33915_1.INJECT1_1 = "NO";
    LUT4 mux_2421_i1_4_lut (.A(n74), .B(n15057[0]), .C(n8478), .D(n52742), 
         .Z(n8479[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i1_4_lut.init = 16'hcfca;
    FD1P3IX pixel_i23 (.D(\Q[10] [23]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[10] [22]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[10] [21]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[10] [20]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[10] [19]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[10] [18]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    FD1P3IX pixel_i17 (.D(\Q[10] [17]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[10] [16]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[10] [15]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[10] [14]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[10] [13]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[10] [12]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[10] [11]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[10] [10]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[10] [9]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[10] [8]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[10] [7]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[10] [6]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[10] [5]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[10] [4]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[10] [3]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[10] [2]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[10] [1]), .SP(sclk_c_enable_2228), .CD(n35688), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2195), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2228), 
            .CD(n35688), .CK(sclk_c), .Q(\RdAddress[10] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_2259), .CD(n35659), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_897), .SP(sclk_c_enable_2259), .CD(n35659), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_2259), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    LUT4 i2433_3_lut (.A(state[2]), .B(state[1]), .C(n13591), .Z(n8478)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2433_3_lut.init = 16'ha8a8;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2410), 
            .CD(n35510), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2410), .CD(n35510), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2410), .CD(n35510), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n8405[4]), .SP(sclk_c_enable_2410), 
            .CD(n35506), .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54979), .SP(sclk_c_enable_2410), .CD(n35506), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=245, LSE_RLINE=245 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    LUT4 mux_2421_i2_4_lut (.A(n71), .B(n15057[0]), .C(n8478), .D(n52742), 
         .Z(n8479[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i2_4_lut.init = 16'hcfca;
    LUT4 mux_2421_i4_4_lut (.A(n38671), .B(n42564), .C(n8478), .D(n4), 
         .Z(n8479[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut_adj_132 (.A(n42702), .B(n54579), .C(n447[3]), .D(n54721), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut_adj_132.init = 16'hfcee;
    LUT4 mux_2421_i8_4_lut (.A(n8303[7]), .B(n42564), .C(n8478), .D(n54579), 
         .Z(n8479[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i8_4_lut.init = 16'h303a;
    LUT4 mux_2421_i9_4_lut (.A(n8303[8]), .B(n42564), .C(n8478), .D(n54579), 
         .Z(n8479[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i9_4_lut.init = 16'h303a;
    LUT4 mux_2421_i10_4_lut (.A(n80), .B(n42564), .C(n8478), .D(n54579), 
         .Z(n8479[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i10_4_lut.init = 16'h303a;
    LUT4 mux_2421_i13_4_lut (.A(n8303[12]), .B(n42564), .C(n8478), .D(n54579), 
         .Z(n8479[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2421_i13_4_lut.init = 16'h303a;
    LUT4 i1_2_lut_rep_617 (.A(state[2]), .B(n13591), .Z(n54620)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_617.init = 16'h4444;
    LUT4 i1_2_lut_rep_576_3_lut (.A(state[2]), .B(n13591), .C(state[1]), 
         .Z(n54579)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_576_3_lut.init = 16'h4040;
    LUT4 i38594_3_lut_rep_582_4_lut (.A(state[2]), .B(n13591), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2410)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38594_3_lut_rep_582_4_lut.init = 16'hfffb;
    PFUMX i38959 (.BLUT(n54977), .ALUT(n54978), .C0(state[1]), .Z(n54979));
    PFUMX i38909 (.BLUT(n54901), .ALUT(n54902), .C0(state[1]), .Z(state_2__N_104[1]));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U35 
//

module \WS2812(48000000,"111111111")_U35  (sclk_c, \port_status[13] , ws2813_out_c_13, 
            state, n54583, \Q[13] , \RdAddress[13] , GND_net);
    input sclk_c;
    output \port_status[13] ;
    output ws2813_out_c_13;
    output [2:0]state;
    input n54583;
    input [23:0]\Q[13] ;
    output [8:0]\RdAddress[13] ;
    input GND_net;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_2125;
    wire [31:0]n9280;
    
    wire sclk_c_enable_121, n54776, sclk_c_enable_122, serial_N_433, 
        sclk_c_enable_126;
    wire [2:0]state_2__N_104;
    wire [31:0]n9104;
    
    wire n42586, n9279, n54592, n53124, n53125;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53128, n53126, n53127, n53129, n13801, n8022;
    wire [31:0]n447;
    
    wire n54845, n13766, n11, n55539;
    wire [6:0]n15081;
    
    wire n55536, n38311, sclk_c_enable_1910;
    wire [31:0]bit_counter_31__N_204;
    wire [31:0]bit_counter_31__N_172;
    
    wire n55535, n54710, n54947, n54946, n54950, n54949, sclk_c_enable_1943, 
        n45, n53, n54844, n53331, n53332, n53333, n1, n52655;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    
    wire n35973;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    wire [8:0]cur_pixel_8__N_107;
    wire [8:0]n118;
    
    wire sclk_c_enable_1974, n47999, n47998, n47997, n47996, n47995, 
        n47994, n47993, n53116, n53117, n53118, n53119, n47992, 
        n53120, n53121, n47991, n1_adj_896, n53122, n53123, n47990, 
        n47989, n47988, n54889, n54890, n47987, n53330, n53329, 
        n53328, n53327, n4, n47986, n47985, n54951, n47984, n53130, 
        serial_N_437, n15, n14, n47634, n47633, n47632, n47631, 
        n35795, n47630, n54948, n54846, n47629, n47628, n47627, 
        n47918, n47917, n47916, n47915, n47626, n47625, n47624, 
        n47623, n47622, n47621, n47620, n47619, n48753, n48752, 
        n48751, n48750, n48749, n48748, n48747, n48746, n48745, 
        n48744, n48743, n48742, n48741, n48740, n48739, n48738, 
        n48689, n48688, n48687, n48686, n48685, n48684, n48683, 
        n48682, n48681, n48680, n48679, n48678, n48677, n48676, 
        n48675, n48674;
    
    FD1P3AX delay_counter_i0_i0 (.D(n9280[0]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54776), .SP(sclk_c_enable_121), .CK(sclk_c), 
            .Q(\port_status[13] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_122), .CK(sclk_c), 
            .Q(ws2813_out_c_13)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_126), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_126), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_126), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    LUT4 mux_2592_i9_4_lut (.A(n9104[8]), .B(n42586), .C(n9279), .D(n54592), 
         .Z(n9280[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i9_4_lut.init = 16'h303a;
    L6MUX21 i37922 (.D0(n53124), .D1(n53125), .SD(bit_counter[2]), .Z(n53128));
    L6MUX21 i37923 (.D0(n53126), .D1(n53127), .SD(bit_counter[2]), .Z(n53129));
    LUT4 i38437_2_lut_3_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .D(n13801), .Z(sclk_c_enable_126)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i38437_2_lut_3_lut_4_lut_4_lut.init = 16'hffc2;
    LUT4 i2345_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n13801), 
         .D(state[0]), .Z(n8022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2345_4_lut_4_lut_4_lut.init = 16'he8c8;
    LUT4 mux_2582_i3_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13801), .Z(n54845)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2582_i3_4_lut_then_4_lut.init = 16'hb1f0;
    LUT4 i1_2_lut_rep_844 (.A(n13766), .B(n11), .Z(n55539)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_844.init = 16'h8888;
    LUT4 i28717_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n15081[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28717_2_lut_3_lut.init = 16'h7070;
    LUT4 i30413_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42586)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i30413_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut_4_lut_then_2_lut (.A(state[2]), .B(n13801), .Z(n55536)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_then_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13766), 
         .D(state[1]), .Z(n38311)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[0]), .B(state[2]), .C(n13766), 
         .D(state[1]), .Z(sclk_c_enable_1910)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'hcc20;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_4_lut_else_2_lut_4_lut (.A(n13766), .B(n11), .C(state[0]), 
         .D(state[2]), .Z(n55535)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_else_2_lut_4_lut.init = 16'h0070;
    LUT4 i1_2_lut_3_lut_adj_55 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_55.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_56 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_56.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_57 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_57.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_58 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_58.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_59 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_59.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_60 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_60.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_61 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_61.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_62 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_62.init = 16'h2020;
    LUT4 mux_2576_i9_3_lut_4_lut (.A(n13766), .B(n11), .C(n54710), .D(n447[8]), 
         .Z(n9104[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2576_i9_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_3_lut_adj_63 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_63.init = 16'h2020;
    LUT4 mux_2576_i10_3_lut_4_lut (.A(n13766), .B(n11), .C(n54710), .D(n447[9]), 
         .Z(n9104[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2576_i10_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_3_lut_adj_64 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_64.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_65 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_65.init = 16'h2020;
    LUT4 mux_2576_i13_3_lut_4_lut (.A(n13766), .B(n11), .C(n54710), .D(n447[12]), 
         .Z(n9104[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_2576_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2582_i5_4_lut_4_lut_then_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13801), .Z(n54947)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2582_i5_4_lut_4_lut_then_4_lut.init = 16'he2e0;
    LUT4 i1_2_lut_3_lut_adj_66 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_66.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_67 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_67.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_68 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_68.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_69 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_69.init = 16'h2020;
    LUT4 mux_2582_i5_4_lut_4_lut_else_4_lut (.A(state[1]), .B(state[2]), 
         .C(n447[4]), .D(n13801), .Z(n54946)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_2582_i5_4_lut_4_lut_else_4_lut.init = 16'hd0f0;
    LUT4 i1_2_lut_3_lut_adj_70 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_70.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_71 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_71.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_72 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_72.init = 16'h2020;
    LUT4 i1_2_lut_rep_589_3_lut (.A(state[2]), .B(n13801), .C(state[1]), 
         .Z(n54592)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_589_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_73.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_then_4_lut (.A(state[2]), .B(state[0]), .C(n447[7]), 
         .D(state[1]), .Z(n54950)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_then_4_lut.init = 16'hf0f4;
    LUT4 i1_3_lut_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[7]), 
         .D(state[1]), .Z(n54949)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_else_4_lut.init = 16'hf0b0;
    LUT4 i1_2_lut_3_lut_adj_74 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_74.init = 16'h2020;
    LUT4 i38587_3_lut_rep_590_4_lut (.A(state[2]), .B(n13801), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_2125)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38587_3_lut_rep_590_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_3_lut_adj_75 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_75.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_76 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_76.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_77 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_77.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_78 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_78.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_79 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_79.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_80 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_80.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_81 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_81.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_82 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_82.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_83 (.A(state[0]), .B(state[2]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_3_lut_adj_83.init = 16'h2020;
    LUT4 i1_2_lut_rep_707_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n54710)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_707_3_lut.init = 16'hefef;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13801), 
         .Z(sclk_c_enable_122)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_3_lut_rep_682_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_1943)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_682_4_lut_3_lut.init = 16'h8989;
    LUT4 i1_2_lut_3_lut_4_lut_adj_84 (.A(state[2]), .B(state[1]), .C(n447[0]), 
         .D(state[0]), .Z(n45)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_84.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_85 (.A(state[2]), .B(state[1]), .C(n447[1]), 
         .D(state[0]), .Z(n53)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_85.init = 16'he0f0;
    LUT4 mux_2582_i3_4_lut_else_4_lut (.A(state[2]), .B(state[0]), .C(n447[2]), 
         .D(n13766), .Z(n54844)) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2582_i3_4_lut_else_4_lut.init = 16'hb0f4;
    LUT4 mux_2592_i10_4_lut (.A(n9104[9]), .B(n42586), .C(n9279), .D(n54592), 
         .Z(n9280[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i10_4_lut.init = 16'h303a;
    L6MUX21 i38127 (.D0(n53331), .D1(n53332), .SD(bit_counter[2]), .Z(n53333));
    LUT4 mux_2338_i2_4_lut_4_lut (.A(n54583), .B(n54710), .C(n8022), .D(n13766), 
         .Z(state_2__N_104[1])) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C)+!B (C+!(D))))) */ ;
    defparam mux_2338_i2_4_lut_4_lut.init = 16'h5053;
    LUT4 i28782_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28782_2_lut.init = 16'hbbbb;
    LUT4 mux_2592_i2_4_lut (.A(n53), .B(n15081[0]), .C(n9279), .D(n52655), 
         .Z(n9280[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i2_4_lut.init = 16'hcfca;
    FD1P3AX delay_counter_i0_i1 (.D(n9280[1]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n9280[3]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n9280[7]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n9280[8]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n9280[9]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n9280[12]), .SP(sclk_c_enable_2125), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3IX pixel_i0 (.D(\Q[13] [0]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    LUT4 i28766_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i28766_2_lut_3_lut.init = 16'h1010;
    LUT4 i29594_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[8]), .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29594_2_lut_3_lut.init = 16'h1010;
    LUT4 i29593_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[7]), .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29593_2_lut_3_lut.init = 16'h1010;
    LUT4 i29605_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[6]), .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29605_2_lut_3_lut.init = 16'h1010;
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    LUT4 i29604_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[5]), .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29604_2_lut_3_lut.init = 16'h1010;
    LUT4 i29639_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[4]), .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29639_2_lut_3_lut.init = 16'h1010;
    LUT4 i29602_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[3]), .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29602_2_lut_3_lut.init = 16'h1010;
    LUT4 i29661_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[2]), .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29661_2_lut_3_lut.init = 16'h1010;
    LUT4 i30126_2_lut_3_lut (.A(state[2]), .B(n11), .C(n118[1]), .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i30126_2_lut_3_lut.init = 16'h1010;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47999), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47998), .COUT(n47999), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47997), .COUT(n47998), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47996), .COUT(n47997), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47995), .COUT(n47996), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47994), .COUT(n47995), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47993), .COUT(n47994), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    PFUMX i37918 (.BLUT(n53116), .ALUT(n53117), .C0(bit_counter[1]), .Z(n53124));
    PFUMX i37919 (.BLUT(n53118), .ALUT(n53119), .C0(bit_counter[1]), .Z(n53125));
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47992), .COUT(n47993), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    PFUMX i37920 (.BLUT(n53120), .ALUT(n53121), .C0(bit_counter[1]), .Z(n53126));
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47991), .COUT(n47992), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    LUT4 i28781_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_896)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28781_2_lut.init = 16'hbbbb;
    PFUMX i37921 (.BLUT(n53122), .ALUT(n53123), .C0(bit_counter[1]), .Z(n53127));
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47990), .COUT(n47991), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47989), .COUT(n47990), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47988), .COUT(n47989), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    PFUMX i38901 (.BLUT(n54889), .ALUT(n54890), .C0(state[1]), .Z(state_2__N_104[2]));
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47987), .COUT(n47988), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    LUT4 i38124_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38124_3_lut.init = 16'hcaca;
    LUT4 i38123_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38123_3_lut.init = 16'hcaca;
    LUT4 i38122_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38122_3_lut.init = 16'hcaca;
    LUT4 i38121_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38121_3_lut.init = 16'hcaca;
    LUT4 mux_2592_i13_4_lut (.A(n9104[12]), .B(n42586), .C(n9279), .D(n54592), 
         .Z(n9280[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i13_4_lut.init = 16'h303a;
    LUT4 mux_2592_i4_4_lut (.A(n38311), .B(n42586), .C(n9279), .D(n4), 
         .Z(n9280[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut (.A(n11), .B(n54592), .C(n447[3]), .D(n54710), .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut.init = 16'hfcee;
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47986), .COUT(n47987), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    LUT4 mux_2338_i3_4_lut_then_3_lut (.A(state[0]), .B(n13801), .C(state[2]), 
         .Z(n54890)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2338_i3_4_lut_then_3_lut.init = 16'h0808;
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47985), .COUT(n47986), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    LUT4 mux_2592_i8_4_lut (.A(n54951), .B(n42586), .C(n9279), .D(n54592), 
         .Z(n9280[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i8_4_lut.init = 16'h303a;
    LUT4 mux_2338_i3_4_lut_else_3_lut (.A(state[0]), .B(state[2]), .C(n11), 
         .D(n13766), .Z(n54889)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2338_i3_4_lut_else_3_lut.init = 16'h2000;
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47984), .COUT(n47985), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47984), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    LUT4 i37917_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37917_3_lut.init = 16'hcaca;
    LUT4 i37916_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37916_3_lut.init = 16'hcaca;
    LUT4 i37915_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37915_3_lut.init = 16'hcaca;
    LUT4 i37914_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37914_3_lut.init = 16'hcaca;
    LUT4 i37913_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37913_3_lut.init = 16'hcaca;
    LUT4 i37912_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37912_3_lut.init = 16'hcaca;
    LUT4 i37911_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37911_3_lut.init = 16'hcaca;
    LUT4 i37910_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37910_3_lut.init = 16'hcaca;
    LUT4 i38408_2_lut_rep_736 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1974)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38408_2_lut_rep_736.init = 16'h9999;
    LUT4 i23732_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35973)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23732_2_lut_2_lut.init = 16'h8888;
    L6MUX21 i37924 (.D0(n53128), .D1(n53129), .SD(bit_counter[3]), .Z(n53130));
    PFUMX i38125 (.BLUT(n53327), .ALUT(n53328), .C0(bit_counter[1]), .Z(n53331));
    PFUMX i38126 (.BLUT(n53329), .ALUT(n53330), .C0(bit_counter[1]), .Z(n53332));
    LUT4 i19533_1_lut_rep_773 (.A(state[2]), .Z(n54776)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i19533_1_lut_rep_773.init = 16'h5555;
    LUT4 i28668_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28668_3_lut_3_lut.init = 16'h5151;
    LUT4 mux_2592_i1_4_lut (.A(n45), .B(n15081[0]), .C(n9279), .D(n52655), 
         .Z(n9280[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2592_i1_4_lut.init = 16'hcfca;
    LUT4 i2604_3_lut (.A(state[2]), .B(state[1]), .C(n13801), .Z(n9279)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i2604_3_lut.init = 16'ha8a8;
    FD1P3IX pixel_i23 (.D(\Q[13] [23]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[13] [22]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    FD1P3IX pixel_i21 (.D(\Q[13] [21]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[13] [20]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[13] [19]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[13] [18]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[8]), .C(n14), .D(cur_pixel[1]), 
         .Z(n11)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    FD1P3IX pixel_i17 (.D(\Q[13] [17]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[13] [16]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    LUT4 i6_4_lut (.A(cur_pixel[0]), .B(cur_pixel[2]), .C(cur_pixel[6]), 
         .D(cur_pixel[7]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    FD1P3IX pixel_i15 (.D(\Q[13] [15]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    LUT4 i5_3_lut (.A(cur_pixel[3]), .B(cur_pixel[5]), .C(cur_pixel[4]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    FD1P3IX pixel_i14 (.D(\Q[13] [14]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[13] [13]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[13] [12]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[13] [11]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[13] [10]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[13] [9]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[13] [8]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[13] [7]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[13] [6]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[13] [5]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[13] [4]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[13] [3]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[13] [2]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[13] [1]), .SP(sclk_c_enable_1943), .CD(n35973), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_1910), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_1943), 
            .CD(n35973), .CK(sclk_c), .Q(\RdAddress[13] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1974), .CD(n35973), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_896), .SP(sclk_c_enable_1974), .CD(n35973), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1974), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    CCU2D add_3128_33 (.A0(bit_counter[31]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47634), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_33.INIT0 = 16'h5999;
    defparam add_3128_33.INIT1 = 16'h0000;
    defparam add_3128_33.INJECT1_0 = "NO";
    defparam add_3128_33.INJECT1_1 = "NO";
    CCU2D add_3128_31 (.A0(bit_counter[29]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47633), .COUT(n47634), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_31.INIT0 = 16'h5999;
    defparam add_3128_31.INIT1 = 16'h5999;
    defparam add_3128_31.INJECT1_0 = "NO";
    defparam add_3128_31.INJECT1_1 = "NO";
    CCU2D add_3128_29 (.A0(bit_counter[27]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47632), .COUT(n47633), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_29.INIT0 = 16'h5999;
    defparam add_3128_29.INIT1 = 16'h5999;
    defparam add_3128_29.INJECT1_0 = "NO";
    defparam add_3128_29.INJECT1_1 = "NO";
    CCU2D add_3128_27 (.A0(bit_counter[25]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47631), .COUT(n47632), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_27.INIT0 = 16'h5999;
    defparam add_3128_27.INIT1 = 16'h5999;
    defparam add_3128_27.INJECT1_0 = "NO";
    defparam add_3128_27.INJECT1_1 = "NO";
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    CCU2D add_3128_25 (.A0(bit_counter[23]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47630), .COUT(n47631), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_25.INIT0 = 16'h5999;
    defparam add_3128_25.INIT1 = 16'h5999;
    defparam add_3128_25.INJECT1_0 = "NO";
    defparam add_3128_25.INJECT1_1 = "NO";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_2125), 
            .CD(n35795), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_2125), .CD(n35795), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_2125), .CD(n35795), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n54948), .SP(sclk_c_enable_2125), .CD(n9279), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54846), .SP(sclk_c_enable_2125), .CD(n9279), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=19, LSE_LLINE=278, LSE_RLINE=278 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    CCU2D add_3128_23 (.A0(bit_counter[21]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47629), .COUT(n47630), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_23.INIT0 = 16'h5999;
    defparam add_3128_23.INIT1 = 16'h5999;
    defparam add_3128_23.INJECT1_0 = "NO";
    defparam add_3128_23.INJECT1_1 = "NO";
    CCU2D add_3128_21 (.A0(bit_counter[19]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47628), .COUT(n47629), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_21.INIT0 = 16'h5999;
    defparam add_3128_21.INIT1 = 16'h5999;
    defparam add_3128_21.INJECT1_0 = "NO";
    defparam add_3128_21.INJECT1_1 = "NO";
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    CCU2D add_3128_19 (.A0(bit_counter[17]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47627), .COUT(n47628), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_19.INIT0 = 16'h5999;
    defparam add_3128_19.INIT1 = 16'h5999;
    defparam add_3128_19.INJECT1_0 = "NO";
    defparam add_3128_19.INJECT1_1 = "NO";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53130), .B(n53333), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47918), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47917), .COUT(n47918), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47916), .COUT(n47917), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47915), .COUT(n47916), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47915), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 mux_2338_i1_4_lut (.A(n54710), .B(n54583), .C(n8022), .D(n55539), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_2338_i1_4_lut.init = 16'h3f3a;
    CCU2D add_3128_17 (.A0(bit_counter[15]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47626), .COUT(n47627), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_17.INIT0 = 16'h5999;
    defparam add_3128_17.INIT1 = 16'h5999;
    defparam add_3128_17.INJECT1_0 = "NO";
    defparam add_3128_17.INJECT1_1 = "NO";
    CCU2D add_3128_15 (.A0(bit_counter[13]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47625), .COUT(n47626), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_15.INIT0 = 16'h5999;
    defparam add_3128_15.INIT1 = 16'h5999;
    defparam add_3128_15.INJECT1_0 = "NO";
    defparam add_3128_15.INJECT1_1 = "NO";
    CCU2D add_3128_13 (.A0(bit_counter[11]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47624), .COUT(n47625), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_13.INIT0 = 16'h5999;
    defparam add_3128_13.INIT1 = 16'h5999;
    defparam add_3128_13.INJECT1_0 = "NO";
    defparam add_3128_13.INJECT1_1 = "NO";
    CCU2D add_3128_11 (.A0(bit_counter[9]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47623), .COUT(n47624), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_11.INIT0 = 16'h5999;
    defparam add_3128_11.INIT1 = 16'h5999;
    defparam add_3128_11.INJECT1_0 = "NO";
    defparam add_3128_11.INJECT1_1 = "NO";
    CCU2D add_3128_9 (.A0(bit_counter[7]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47622), .COUT(n47623), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_9.INIT0 = 16'h5999;
    defparam add_3128_9.INIT1 = 16'h5999;
    defparam add_3128_9.INJECT1_0 = "NO";
    defparam add_3128_9.INJECT1_1 = "NO";
    CCU2D add_3128_7 (.A0(bit_counter[5]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47621), .COUT(n47622), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_7.INIT0 = 16'h5999;
    defparam add_3128_7.INIT1 = 16'h5999;
    defparam add_3128_7.INJECT1_0 = "NO";
    defparam add_3128_7.INJECT1_1 = "NO";
    CCU2D add_3128_5 (.A0(bit_counter[3]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47620), .COUT(n47621), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_5.INIT0 = 16'h5999;
    defparam add_3128_5.INIT1 = 16'h5999;
    defparam add_3128_5.INJECT1_0 = "NO";
    defparam add_3128_5.INJECT1_1 = "NO";
    CCU2D add_3128_3 (.A0(bit_counter[1]), .B0(n13766), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13766), .C1(GND_net), 
          .D1(GND_net), .CIN(n47619), .COUT(n47620), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_3.INIT0 = 16'h5999;
    defparam add_3128_3.INIT1 = 16'h5999;
    defparam add_3128_3.INJECT1_0 = "NO";
    defparam add_3128_3.INJECT1_1 = "NO";
    CCU2D add_3128_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13766), .C1(GND_net), .D1(GND_net), 
          .COUT(n47619), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3128_1.INIT0 = 16'hF000;
    defparam add_3128_1.INIT1 = 16'h5999;
    defparam add_3128_1.INJECT1_0 = "NO";
    defparam add_3128_1.INJECT1_1 = "NO";
    PFUMX i38871 (.BLUT(n54844), .ALUT(n54845), .C0(state[1]), .Z(n54846));
    CCU2D add_33906_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48753), 
          .S0(n13801));
    defparam add_33906_cout.INIT0 = 16'h0000;
    defparam add_33906_cout.INIT1 = 16'h0000;
    defparam add_33906_cout.INJECT1_0 = "NO";
    defparam add_33906_cout.INJECT1_1 = "NO";
    CCU2D add_33906_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48752), .COUT(n48753));
    defparam add_33906_31.INIT0 = 16'hf555;
    defparam add_33906_31.INIT1 = 16'h5555;
    defparam add_33906_31.INJECT1_0 = "NO";
    defparam add_33906_31.INJECT1_1 = "NO";
    CCU2D add_33906_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48751), .COUT(n48752));
    defparam add_33906_29.INIT0 = 16'hf555;
    defparam add_33906_29.INIT1 = 16'hf555;
    defparam add_33906_29.INJECT1_0 = "NO";
    defparam add_33906_29.INJECT1_1 = "NO";
    CCU2D add_33906_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48750), .COUT(n48751));
    defparam add_33906_27.INIT0 = 16'hf555;
    defparam add_33906_27.INIT1 = 16'hf555;
    defparam add_33906_27.INJECT1_0 = "NO";
    defparam add_33906_27.INJECT1_1 = "NO";
    CCU2D add_33906_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48749), .COUT(n48750));
    defparam add_33906_25.INIT0 = 16'hf555;
    defparam add_33906_25.INIT1 = 16'hf555;
    defparam add_33906_25.INJECT1_0 = "NO";
    defparam add_33906_25.INJECT1_1 = "NO";
    CCU2D add_33906_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48748), .COUT(n48749));
    defparam add_33906_23.INIT0 = 16'hf555;
    defparam add_33906_23.INIT1 = 16'hf555;
    defparam add_33906_23.INJECT1_0 = "NO";
    defparam add_33906_23.INJECT1_1 = "NO";
    CCU2D add_33906_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48747), .COUT(n48748));
    defparam add_33906_21.INIT0 = 16'hf555;
    defparam add_33906_21.INIT1 = 16'hf555;
    defparam add_33906_21.INJECT1_0 = "NO";
    defparam add_33906_21.INJECT1_1 = "NO";
    CCU2D add_33906_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48746), .COUT(n48747));
    defparam add_33906_19.INIT0 = 16'hf555;
    defparam add_33906_19.INIT1 = 16'hf555;
    defparam add_33906_19.INJECT1_0 = "NO";
    defparam add_33906_19.INJECT1_1 = "NO";
    CCU2D add_33906_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48745), .COUT(n48746));
    defparam add_33906_17.INIT0 = 16'hf555;
    defparam add_33906_17.INIT1 = 16'hf555;
    defparam add_33906_17.INJECT1_0 = "NO";
    defparam add_33906_17.INJECT1_1 = "NO";
    CCU2D add_33906_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48744), .COUT(n48745));
    defparam add_33906_15.INIT0 = 16'hf555;
    defparam add_33906_15.INIT1 = 16'hf555;
    defparam add_33906_15.INJECT1_0 = "NO";
    defparam add_33906_15.INJECT1_1 = "NO";
    CCU2D add_33906_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48743), .COUT(n48744));
    defparam add_33906_13.INIT0 = 16'hf555;
    defparam add_33906_13.INIT1 = 16'hf555;
    defparam add_33906_13.INJECT1_0 = "NO";
    defparam add_33906_13.INJECT1_1 = "NO";
    CCU2D add_33906_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48742), .COUT(n48743));
    defparam add_33906_11.INIT0 = 16'hf555;
    defparam add_33906_11.INIT1 = 16'hf555;
    defparam add_33906_11.INJECT1_0 = "NO";
    defparam add_33906_11.INJECT1_1 = "NO";
    CCU2D add_33906_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48741), .COUT(n48742));
    defparam add_33906_9.INIT0 = 16'hf555;
    defparam add_33906_9.INIT1 = 16'hf555;
    defparam add_33906_9.INJECT1_0 = "NO";
    defparam add_33906_9.INJECT1_1 = "NO";
    CCU2D add_33906_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48740), .COUT(n48741));
    defparam add_33906_7.INIT0 = 16'hf555;
    defparam add_33906_7.INIT1 = 16'hf555;
    defparam add_33906_7.INJECT1_0 = "NO";
    defparam add_33906_7.INJECT1_1 = "NO";
    CCU2D add_33906_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48739), .COUT(n48740));
    defparam add_33906_5.INIT0 = 16'hf555;
    defparam add_33906_5.INIT1 = 16'hf555;
    defparam add_33906_5.INJECT1_0 = "NO";
    defparam add_33906_5.INJECT1_1 = "NO";
    CCU2D add_33906_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48738), .COUT(n48739));
    defparam add_33906_3.INIT0 = 16'hf555;
    defparam add_33906_3.INIT1 = 16'hf555;
    defparam add_33906_3.INJECT1_0 = "NO";
    defparam add_33906_3.INJECT1_1 = "NO";
    CCU2D add_33906_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n48738));
    defparam add_33906_1.INIT0 = 16'hF000;
    defparam add_33906_1.INIT1 = 16'ha666;
    defparam add_33906_1.INJECT1_0 = "NO";
    defparam add_33906_1.INJECT1_1 = "NO";
    CCU2D add_33907_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n48689), 
          .S0(n13766));
    defparam add_33907_cout.INIT0 = 16'h0000;
    defparam add_33907_cout.INIT1 = 16'h0000;
    defparam add_33907_cout.INJECT1_0 = "NO";
    defparam add_33907_cout.INJECT1_1 = "NO";
    CCU2D add_33907_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48688), .COUT(n48689));
    defparam add_33907_31.INIT0 = 16'hf555;
    defparam add_33907_31.INIT1 = 16'h5555;
    defparam add_33907_31.INJECT1_0 = "NO";
    defparam add_33907_31.INJECT1_1 = "NO";
    CCU2D add_33907_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48687), .COUT(n48688));
    defparam add_33907_29.INIT0 = 16'hf555;
    defparam add_33907_29.INIT1 = 16'hf555;
    defparam add_33907_29.INJECT1_0 = "NO";
    defparam add_33907_29.INJECT1_1 = "NO";
    CCU2D add_33907_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48686), .COUT(n48687));
    defparam add_33907_27.INIT0 = 16'hf555;
    defparam add_33907_27.INIT1 = 16'hf555;
    defparam add_33907_27.INJECT1_0 = "NO";
    defparam add_33907_27.INJECT1_1 = "NO";
    CCU2D add_33907_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48685), .COUT(n48686));
    defparam add_33907_25.INIT0 = 16'hf555;
    defparam add_33907_25.INIT1 = 16'hf555;
    defparam add_33907_25.INJECT1_0 = "NO";
    defparam add_33907_25.INJECT1_1 = "NO";
    CCU2D add_33907_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48684), .COUT(n48685));
    defparam add_33907_23.INIT0 = 16'hf555;
    defparam add_33907_23.INIT1 = 16'hf555;
    defparam add_33907_23.INJECT1_0 = "NO";
    defparam add_33907_23.INJECT1_1 = "NO";
    CCU2D add_33907_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48683), .COUT(n48684));
    defparam add_33907_21.INIT0 = 16'hf555;
    defparam add_33907_21.INIT1 = 16'hf555;
    defparam add_33907_21.INJECT1_0 = "NO";
    defparam add_33907_21.INJECT1_1 = "NO";
    CCU2D add_33907_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48682), .COUT(n48683));
    defparam add_33907_19.INIT0 = 16'hf555;
    defparam add_33907_19.INIT1 = 16'hf555;
    defparam add_33907_19.INJECT1_0 = "NO";
    defparam add_33907_19.INJECT1_1 = "NO";
    CCU2D add_33907_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48681), .COUT(n48682));
    defparam add_33907_17.INIT0 = 16'hf555;
    defparam add_33907_17.INIT1 = 16'hf555;
    defparam add_33907_17.INJECT1_0 = "NO";
    defparam add_33907_17.INJECT1_1 = "NO";
    CCU2D add_33907_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48680), .COUT(n48681));
    defparam add_33907_15.INIT0 = 16'hf555;
    defparam add_33907_15.INIT1 = 16'hf555;
    defparam add_33907_15.INJECT1_0 = "NO";
    defparam add_33907_15.INJECT1_1 = "NO";
    CCU2D add_33907_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48679), .COUT(n48680));
    defparam add_33907_13.INIT0 = 16'hf555;
    defparam add_33907_13.INIT1 = 16'hf555;
    defparam add_33907_13.INJECT1_0 = "NO";
    defparam add_33907_13.INJECT1_1 = "NO";
    CCU2D add_33907_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48678), .COUT(n48679));
    defparam add_33907_11.INIT0 = 16'hf555;
    defparam add_33907_11.INIT1 = 16'hf555;
    defparam add_33907_11.INJECT1_0 = "NO";
    defparam add_33907_11.INJECT1_1 = "NO";
    CCU2D add_33907_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48677), .COUT(n48678));
    defparam add_33907_9.INIT0 = 16'hf555;
    defparam add_33907_9.INIT1 = 16'hf555;
    defparam add_33907_9.INJECT1_0 = "NO";
    defparam add_33907_9.INJECT1_1 = "NO";
    CCU2D add_33907_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48676), .COUT(n48677));
    defparam add_33907_7.INIT0 = 16'hf555;
    defparam add_33907_7.INIT1 = 16'hf555;
    defparam add_33907_7.INJECT1_0 = "NO";
    defparam add_33907_7.INJECT1_1 = "NO";
    CCU2D add_33907_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48675), .COUT(n48676));
    defparam add_33907_5.INIT0 = 16'hf555;
    defparam add_33907_5.INIT1 = 16'hf555;
    defparam add_33907_5.INJECT1_0 = "NO";
    defparam add_33907_5.INJECT1_1 = "NO";
    CCU2D add_33907_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n48674), .COUT(n48675));
    defparam add_33907_3.INIT0 = 16'hf555;
    defparam add_33907_3.INIT1 = 16'hf555;
    defparam add_33907_3.INJECT1_0 = "NO";
    defparam add_33907_3.INJECT1_1 = "NO";
    CCU2D add_33907_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n48674));
    defparam add_33907_1.INIT0 = 16'hF000;
    defparam add_33907_1.INIT1 = 16'ha666;
    defparam add_33907_1.INJECT1_0 = "NO";
    defparam add_33907_1.INJECT1_1 = "NO";
    LUT4 i23603_4_lut (.A(sclk_c_enable_2125), .B(n54592), .C(n9279), 
         .D(n54710), .Z(n35795)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23603_4_lut.init = 16'ha8aa;
    PFUMX i38941 (.BLUT(n54949), .ALUT(n54950), .C0(n55539), .Z(n54951));
    PFUMX i38939 (.BLUT(n54946), .ALUT(n54947), .C0(state[0]), .Z(n54948));
    PFUMX i39243 (.BLUT(n55535), .ALUT(n55536), .C0(state[1]), .Z(n52655));
    
endmodule
//
// Verilog Description of module \WS2812(48000000,"111111111")_U21 
//

module \WS2812(48000000,"111111111")_U21  (\RdAddress[7] , sclk_c, \port_status[7] , 
            ws2813_out_c_7, GND_net, \Q[7] );
    output [8:0]\RdAddress[7] ;
    input sclk_c;
    output \port_status[7] ;
    output ws2813_out_c_7;
    input GND_net;
    input [23:0]\Q[7] ;
    
    wire sclk_c /* synthesis is_clock=1, SET_AS_NETWORK=sclk_c */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/main.vhd(8[3:7])
    
    wire sclk_c_enable_2472, n35403;
    wire [8:0]cur_pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(43[12:21])
    
    wire n53034, n53035;
    wire [31:0]bit_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(46[12:23])
    
    wire n53038, sclk_c_enable_1182;
    wire [31:0]bit_counter_31__N_172;
    wire [31:0]delay_counter;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(45[12:25])
    
    wire sclk_c_enable_960;
    wire [31:0]n6298;
    
    wire sclk_c_enable_70, n54796, sclk_c_enable_71, serial_N_433;
    wire [2:0]state;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    
    wire sclk_c_enable_74;
    wire [2:0]state_2__N_104;
    
    wire n53036, n53037, n53039, n1, n1_adj_895, n48290, n13346;
    wire [31:0]bit_counter_31__N_204;
    
    wire n48289, n48288, n48287, n48286, n48285, n48284, n48283, 
        n48282, n13381, n48281, n48280, sclk_c_enable_2480, n48279, 
        n48278, n48277, n54908, n54907, n54651, n54747, n54663, 
        n35225;
    wire [31:0]n447;
    
    wire n54984, n54983, serial_N_437, n42806, n53289, n53290, n53291, 
        n54595, n54664, n48276, n54609, n35221;
    wire [31:0]n6224;
    
    wire n54985, n48275, n54725;
    wire [31:0]n6122;
    
    wire n80;
    wire [23:0]pixel;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(44[12:17])
    wire [8:0]cur_pixel_8__N_107;
    
    wire n53026, n53027, n53028, n53029, n53030, n53031, n53032, 
        n53033;
    wire [8:0]n118;
    
    wire n54839, n71, n6297, n74;
    wire [6:0]n14750;
    
    wire n42478, n52736, n15, n14, n53288, n53287, n53286, n53285;
    wire [2:0]n9385;
    
    wire n53040, n49102, n49101, n49100, n49099, n49098, n49097, 
        n49096, n49095, n49094, n49093, n49092, n49091, n49090, 
        n49089, n49088, n49087, n49086, n49085, n49084, n49083, 
        n49082, n49081, n49080, n49079, n49078, n39073, n49077, 
        n49076, n49075, n9392, n49074, n49073, n49072, n49071, 
        n47729, n47728, n47727, n47726, n47725, n47724, n47723, 
        n47722, n47721, n47720, n47719, n47718, n47717, n47716, 
        n47715, n47714, n47712, n47711, n4, n47710, n47709;
    
    FD1P3IX PixelAddress_i8 (.D(cur_pixel[8]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [8])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i8.GSR = "DISABLED";
    FD1P3IX PixelAddress_i7 (.D(cur_pixel[7]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [7])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i7.GSR = "DISABLED";
    FD1P3IX PixelAddress_i6 (.D(cur_pixel[6]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [6])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i6.GSR = "DISABLED";
    FD1P3IX PixelAddress_i5 (.D(cur_pixel[5]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i5.GSR = "DISABLED";
    FD1P3IX PixelAddress_i4 (.D(cur_pixel[4]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i4.GSR = "DISABLED";
    FD1P3IX PixelAddress_i3 (.D(cur_pixel[3]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i3.GSR = "DISABLED";
    L6MUX21 i37832 (.D0(n53034), .D1(n53035), .SD(bit_counter[2]), .Z(n53038));
    FD1P3IX PixelAddress_i2 (.D(cur_pixel[2]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i2.GSR = "DISABLED";
    FD1P3IX PixelAddress_i1 (.D(cur_pixel[1]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i1.GSR = "DISABLED";
    FD1P3AX bit_counter_i31 (.D(bit_counter_31__N_172[31]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i31.GSR = "DISABLED";
    FD1P3AX bit_counter_i30 (.D(bit_counter_31__N_172[30]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i30.GSR = "DISABLED";
    FD1P3AX bit_counter_i29 (.D(bit_counter_31__N_172[29]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i29.GSR = "DISABLED";
    FD1P3AX bit_counter_i28 (.D(bit_counter_31__N_172[28]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i28.GSR = "DISABLED";
    FD1P3AX bit_counter_i27 (.D(bit_counter_31__N_172[27]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i27.GSR = "DISABLED";
    FD1P3AX bit_counter_i26 (.D(bit_counter_31__N_172[26]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i26.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i0 (.D(n6298[0]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i25 (.D(bit_counter_31__N_172[25]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i25.GSR = "DISABLED";
    FD1P3AX bit_counter_i24 (.D(bit_counter_31__N_172[24]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i24.GSR = "DISABLED";
    FD1P3AX bit_counter_i23 (.D(bit_counter_31__N_172[23]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i23.GSR = "DISABLED";
    FD1P3AX bit_counter_i22 (.D(bit_counter_31__N_172[22]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i22.GSR = "DISABLED";
    FD1P3AX bit_counter_i21 (.D(bit_counter_31__N_172[21]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i21.GSR = "DISABLED";
    FD1P3AX bit_counter_i20 (.D(bit_counter_31__N_172[20]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i20.GSR = "DISABLED";
    FD1P3AX status_77 (.D(n54796), .SP(sclk_c_enable_70), .CK(sclk_c), 
            .Q(\port_status[7] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam status_77.GSR = "DISABLED";
    FD1P3AX serial_79 (.D(serial_N_433), .SP(sclk_c_enable_71), .CK(sclk_c), 
            .Q(ws2813_out_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam serial_79.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_2__N_104[0]), .SP(sclk_c_enable_74), .CK(sclk_c), 
            .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i0.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(state_2__N_104[1]), .SP(sclk_c_enable_74), .CK(sclk_c), 
            .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_2__N_104[2]), .SP(sclk_c_enable_74), .CK(sclk_c), 
            .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i19 (.D(bit_counter_31__N_172[19]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i19.GSR = "DISABLED";
    L6MUX21 i37833 (.D0(n53036), .D1(n53037), .SD(bit_counter[2]), .Z(n53039));
    FD1P3AX bit_counter_i18 (.D(bit_counter_31__N_172[18]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i18.GSR = "DISABLED";
    FD1P3AX bit_counter_i17 (.D(bit_counter_31__N_172[17]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i17.GSR = "DISABLED";
    FD1P3AX bit_counter_i16 (.D(bit_counter_31__N_172[16]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i16.GSR = "DISABLED";
    FD1P3AX bit_counter_i15 (.D(bit_counter_31__N_172[15]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i15.GSR = "DISABLED";
    FD1P3AX bit_counter_i14 (.D(bit_counter_31__N_172[14]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i14.GSR = "DISABLED";
    FD1P3AX bit_counter_i13 (.D(bit_counter_31__N_172[13]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i13.GSR = "DISABLED";
    FD1P3AX bit_counter_i12 (.D(bit_counter_31__N_172[12]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i12.GSR = "DISABLED";
    FD1P3AX bit_counter_i11 (.D(bit_counter_31__N_172[11]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i11.GSR = "DISABLED";
    FD1P3AX bit_counter_i10 (.D(bit_counter_31__N_172[10]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i10.GSR = "DISABLED";
    FD1P3AX bit_counter_i9 (.D(bit_counter_31__N_172[9]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i9.GSR = "DISABLED";
    FD1P3AX bit_counter_i8 (.D(bit_counter_31__N_172[8]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i8.GSR = "DISABLED";
    FD1P3AX bit_counter_i7 (.D(bit_counter_31__N_172[7]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i7.GSR = "DISABLED";
    FD1P3AX bit_counter_i6 (.D(bit_counter_31__N_172[6]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i6.GSR = "DISABLED";
    FD1P3AX bit_counter_i5 (.D(bit_counter_31__N_172[5]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i5.GSR = "DISABLED";
    FD1P3IX bit_counter_i4 (.D(n1), .SP(sclk_c_enable_1182), .CD(n35403), 
            .CK(sclk_c), .Q(bit_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i4.GSR = "DISABLED";
    FD1P3IX bit_counter_i3 (.D(n1_adj_895), .SP(sclk_c_enable_1182), .CD(n35403), 
            .CK(sclk_c), .Q(bit_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i3.GSR = "DISABLED";
    FD1P3AX bit_counter_i2 (.D(bit_counter_31__N_172[2]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i2.GSR = "DISABLED";
    FD1P3AX bit_counter_i1 (.D(bit_counter_31__N_172[1]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i1.GSR = "DISABLED";
    CCU2D add_3116_33 (.A0(bit_counter[31]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n48290), .S0(bit_counter_31__N_204[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_33.INIT0 = 16'h5999;
    defparam add_3116_33.INIT1 = 16'h0000;
    defparam add_3116_33.INJECT1_0 = "NO";
    defparam add_3116_33.INJECT1_1 = "NO";
    CCU2D add_3116_31 (.A0(bit_counter[29]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[30]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48289), .COUT(n48290), .S0(bit_counter_31__N_204[29]), 
          .S1(bit_counter_31__N_204[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_31.INIT0 = 16'h5999;
    defparam add_3116_31.INIT1 = 16'h5999;
    defparam add_3116_31.INJECT1_0 = "NO";
    defparam add_3116_31.INJECT1_1 = "NO";
    CCU2D add_3116_29 (.A0(bit_counter[27]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[28]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48288), .COUT(n48289), .S0(bit_counter_31__N_204[27]), 
          .S1(bit_counter_31__N_204[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_29.INIT0 = 16'h5999;
    defparam add_3116_29.INIT1 = 16'h5999;
    defparam add_3116_29.INJECT1_0 = "NO";
    defparam add_3116_29.INJECT1_1 = "NO";
    CCU2D add_3116_27 (.A0(bit_counter[25]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[26]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48287), .COUT(n48288), .S0(bit_counter_31__N_204[25]), 
          .S1(bit_counter_31__N_204[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_27.INIT0 = 16'h5999;
    defparam add_3116_27.INIT1 = 16'h5999;
    defparam add_3116_27.INJECT1_0 = "NO";
    defparam add_3116_27.INJECT1_1 = "NO";
    CCU2D add_3116_25 (.A0(bit_counter[23]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[24]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48286), .COUT(n48287), .S0(bit_counter_31__N_204[23]), 
          .S1(bit_counter_31__N_204[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_25.INIT0 = 16'h5999;
    defparam add_3116_25.INIT1 = 16'h5999;
    defparam add_3116_25.INJECT1_0 = "NO";
    defparam add_3116_25.INJECT1_1 = "NO";
    CCU2D add_3116_23 (.A0(bit_counter[21]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[22]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48285), .COUT(n48286), .S0(bit_counter_31__N_204[21]), 
          .S1(bit_counter_31__N_204[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_23.INIT0 = 16'h5999;
    defparam add_3116_23.INIT1 = 16'h5999;
    defparam add_3116_23.INJECT1_0 = "NO";
    defparam add_3116_23.INJECT1_1 = "NO";
    CCU2D add_3116_21 (.A0(bit_counter[19]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[20]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48284), .COUT(n48285), .S0(bit_counter_31__N_204[19]), 
          .S1(bit_counter_31__N_204[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_21.INIT0 = 16'h5999;
    defparam add_3116_21.INIT1 = 16'h5999;
    defparam add_3116_21.INJECT1_0 = "NO";
    defparam add_3116_21.INJECT1_1 = "NO";
    CCU2D add_3116_19 (.A0(bit_counter[17]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[18]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48283), .COUT(n48284), .S0(bit_counter_31__N_204[17]), 
          .S1(bit_counter_31__N_204[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_19.INIT0 = 16'h5999;
    defparam add_3116_19.INIT1 = 16'h5999;
    defparam add_3116_19.INJECT1_0 = "NO";
    defparam add_3116_19.INJECT1_1 = "NO";
    CCU2D add_3116_17 (.A0(bit_counter[15]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[16]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48282), .COUT(n48283), .S0(bit_counter_31__N_204[15]), 
          .S1(bit_counter_31__N_204[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_17.INIT0 = 16'h5999;
    defparam add_3116_17.INIT1 = 16'h5999;
    defparam add_3116_17.INJECT1_0 = "NO";
    defparam add_3116_17.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .D(n13381), .Z(sclk_c_enable_74)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hffc2;
    CCU2D add_3116_15 (.A0(bit_counter[13]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[14]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48281), .COUT(n48282), .S0(bit_counter_31__N_204[13]), 
          .S1(bit_counter_31__N_204[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_15.INIT0 = 16'h5999;
    defparam add_3116_15.INIT1 = 16'h5999;
    defparam add_3116_15.INJECT1_0 = "NO";
    defparam add_3116_15.INJECT1_1 = "NO";
    CCU2D add_3116_13 (.A0(bit_counter[11]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[12]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48280), .COUT(n48281), .S0(bit_counter_31__N_204[11]), 
          .S1(bit_counter_31__N_204[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_13.INIT0 = 16'h5999;
    defparam add_3116_13.INIT1 = 16'h5999;
    defparam add_3116_13.INJECT1_0 = "NO";
    defparam add_3116_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(n13346), 
         .D(state[0]), .Z(sclk_c_enable_2480)) /* synthesis lut_function=(A (B)+!A !(B+!(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h9888;
    CCU2D add_3116_11 (.A0(bit_counter[9]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[10]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48279), .COUT(n48280), .S0(bit_counter_31__N_204[9]), 
          .S1(bit_counter_31__N_204[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_11.INIT0 = 16'h5999;
    defparam add_3116_11.INIT1 = 16'h5999;
    defparam add_3116_11.INJECT1_0 = "NO";
    defparam add_3116_11.INJECT1_1 = "NO";
    CCU2D add_3116_9 (.A0(bit_counter[7]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[8]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48278), .COUT(n48279), .S0(bit_counter_31__N_204[7]), 
          .S1(bit_counter_31__N_204[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_9.INIT0 = 16'h5999;
    defparam add_3116_9.INIT1 = 16'h5999;
    defparam add_3116_9.INJECT1_0 = "NO";
    defparam add_3116_9.INJECT1_1 = "NO";
    CCU2D add_3116_7 (.A0(bit_counter[5]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[6]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48277), .COUT(n48278), .S0(bit_counter_31__N_204[5]), 
          .S1(bit_counter_31__N_204[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_7.INIT0 = 16'h5999;
    defparam add_3116_7.INIT1 = 16'h5999;
    defparam add_3116_7.INJECT1_0 = "NO";
    defparam add_3116_7.INJECT1_1 = "NO";
    LUT4 i38583_4_lut_then_3_lut (.A(state[2]), .B(state[0]), .C(n13381), 
         .Z(n54908)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i38583_4_lut_then_3_lut.init = 16'h1010;
    LUT4 i38583_4_lut_else_3_lut (.A(state[2]), .B(state[0]), .C(n13346), 
         .Z(n54907)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i38583_4_lut_else_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_648 (.A(state[1]), .B(n13381), .Z(n54651)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_648.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[1]), .B(n13381), .C(n54747), .D(n54663), 
         .Z(state_2__N_104[2])) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd080;
    FD1P3IX delay_counter_i0_i31 (.D(n447[31]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i31.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i30 (.D(n447[30]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i30.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i29 (.D(n447[29]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i29.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i28 (.D(n447[28]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i28.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i27 (.D(n447[27]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i27.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i26 (.D(n447[26]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i26.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i25 (.D(n447[25]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i25.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i24 (.D(n447[24]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i24.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i23 (.D(n447[23]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i23.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i22 (.D(n447[22]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i22.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i21 (.D(n447[21]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i21.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i20 (.D(n447[20]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i20.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i19 (.D(n447[19]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i19.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i18 (.D(n447[18]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i18.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i17 (.D(n447[17]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i17.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i16 (.D(n447[16]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i16.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i15 (.D(n447[15]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i15.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i14 (.D(n447[14]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i14.GSR = "DISABLED";
    LUT4 mux_1928_i3_4_lut_then_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13381), .Z(n54984)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1928_i3_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 mux_1928_i3_4_lut_else_4_lut (.A(state[0]), .B(state[2]), .C(n447[2]), 
         .D(n13346), .Z(n54983)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1928_i3_4_lut_else_4_lut.init = 16'hd0f2;
    FD1P3IX delay_counter_i0_i13 (.D(n447[13]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i13.GSR = "DISABLED";
    LUT4 i26876_1_lut_rep_793 (.A(state[2]), .Z(n54796)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i26876_1_lut_rep_793.init = 16'h5555;
    LUT4 i28919_3_lut_3_lut (.A(state[2]), .B(state[0]), .C(serial_N_437), 
         .Z(serial_N_433)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i28919_3_lut_3_lut.init = 16'h5151;
    LUT4 i1_2_lut_rep_660 (.A(n42806), .B(n13346), .Z(n54663)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_660.init = 16'h8888;
    L6MUX21 i38085 (.D0(n53289), .D1(n53290), .SD(bit_counter[2]), .Z(n53291));
    LUT4 i1_2_lut_rep_592_3_lut (.A(n42806), .B(n13346), .C(state[1]), 
         .Z(n54595)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_592_3_lut.init = 16'h0808;
    FD1P3IX delay_counter_i0_i11 (.D(n447[11]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i11.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_661 (.A(state[2]), .B(n13381), .Z(n54664)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_661.init = 16'h4444;
    CCU2D add_3116_5 (.A0(bit_counter[3]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[4]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48276), .COUT(n48277), .S0(bit_counter_31__N_204[3]), 
          .S1(bit_counter_31__N_204[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_5.INIT0 = 16'h5999;
    defparam add_3116_5.INIT1 = 16'h5999;
    defparam add_3116_5.INJECT1_0 = "NO";
    defparam add_3116_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_606_3_lut (.A(state[2]), .B(n13381), .C(state[1]), 
         .Z(n54609)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_2_lut_rep_606_3_lut.init = 16'h4040;
    FD1P3IX delay_counter_i0_i10 (.D(n447[10]), .SP(sclk_c_enable_960), 
            .CD(n35225), .CK(sclk_c), .Q(delay_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i10.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i6 (.D(n447[6]), .SP(sclk_c_enable_960), .CD(n35225), 
            .CK(sclk_c), .Q(delay_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i6.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i5 (.D(n447[5]), .SP(sclk_c_enable_960), .CD(n35225), 
            .CK(sclk_c), .Q(delay_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i5.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i4 (.D(n6224[4]), .SP(sclk_c_enable_960), .CD(n35221), 
            .CK(sclk_c), .Q(delay_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i4.GSR = "DISABLED";
    FD1P3IX delay_counter_i0_i2 (.D(n54985), .SP(sclk_c_enable_960), .CD(n35221), 
            .CK(sclk_c), .Q(delay_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i2.GSR = "DISABLED";
    CCU2D add_3116_3 (.A0(bit_counter[1]), .B0(n13346), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[2]), .B1(n13346), .C1(GND_net), 
          .D1(GND_net), .CIN(n48275), .COUT(n48276), .S0(bit_counter_31__N_204[1]), 
          .S1(bit_counter_31__N_204[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_3.INIT0 = 16'h5999;
    defparam add_3116_3.INIT1 = 16'h5999;
    defparam add_3116_3.INJECT1_0 = "NO";
    defparam add_3116_3.INJECT1_1 = "NO";
    LUT4 i38600_3_lut_rep_607_4_lut (.A(state[2]), .B(n13381), .C(state[1]), 
         .D(state[0]), .Z(sclk_c_enable_960)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i38600_3_lut_rep_607_4_lut.init = 16'hfffb;
    CCU2D add_3116_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(n13346), .C1(GND_net), .D1(GND_net), 
          .COUT(n48275), .S1(bit_counter_31__N_204[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(63[5] 77[12])
    defparam add_3116_1.INIT0 = 16'hF000;
    defparam add_3116_1.INIT1 = 16'h5999;
    defparam add_3116_1.INJECT1_0 = "NO";
    defparam add_3116_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(n54595), .B(n54747), .C(n447[8]), .D(n54725), 
         .Z(n6122[8])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_8 (.A(n54595), .B(n54747), .C(n447[12]), .D(n54725), 
         .Z(n6122[12])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_8.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_9 (.A(n54595), .B(n54747), .C(n447[9]), .D(n54725), 
         .Z(n80)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_9.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_10 (.A(n54595), .B(n54747), .C(n447[7]), .D(n54725), 
         .Z(n6122[7])) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_adj_10.init = 16'hf888;
    FD1P3AX delay_counter_i0_i1 (.D(n6298[1]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i1.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i3 (.D(n6298[3]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i3.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i7 (.D(n6298[7]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i7.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i8 (.D(n6298[8]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i8.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i9 (.D(n6298[9]), .SP(sclk_c_enable_960), .CK(sclk_c), 
            .Q(delay_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i9.GSR = "DISABLED";
    FD1P3AX delay_counter_i0_i12 (.D(n6298[12]), .SP(sclk_c_enable_960), 
            .CK(sclk_c), .Q(delay_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam delay_counter_i0_i12.GSR = "DISABLED";
    FD1P3IX pixel_i0 (.D(\Q[7] [0]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i0.GSR = "DISABLED";
    FD1P3AX cur_pixel_i0 (.D(cur_pixel_8__N_107[0]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i0.GSR = "DISABLED";
    FD1P3IX PixelAddress_i0 (.D(cur_pixel[0]), .SP(sclk_c_enable_2472), 
            .CD(n35403), .CK(sclk_c), .Q(\RdAddress[7] [0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam PixelAddress_i0.GSR = "DISABLED";
    FD1P3AX bit_counter_i0 (.D(bit_counter_31__N_172[0]), .SP(sclk_c_enable_1182), 
            .CK(sclk_c), .Q(bit_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam bit_counter_i0.GSR = "DISABLED";
    PFUMX i37828 (.BLUT(n53026), .ALUT(n53027), .C0(bit_counter[1]), .Z(n53034));
    PFUMX i37829 (.BLUT(n53028), .ALUT(n53029), .C0(bit_counter[1]), .Z(n53035));
    PFUMX i37830 (.BLUT(n53030), .ALUT(n53031), .C0(bit_counter[1]), .Z(n53036));
    PFUMX i37831 (.BLUT(n53032), .ALUT(n53033), .C0(bit_counter[1]), .Z(n53037));
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n42806), .C(n118[0]), .Z(cur_pixel_8__N_107[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_11 (.A(state[2]), .B(n42806), .C(n118[8]), 
         .Z(cur_pixel_8__N_107[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_11.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_12 (.A(state[2]), .B(n42806), .C(n118[7]), 
         .Z(cur_pixel_8__N_107[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_12.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_13 (.A(state[2]), .B(n42806), .C(n118[6]), 
         .Z(cur_pixel_8__N_107[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_13.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_14 (.A(state[2]), .B(n42806), .C(n118[5]), 
         .Z(cur_pixel_8__N_107[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_14.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_15 (.A(state[2]), .B(n42806), .C(n118[4]), 
         .Z(cur_pixel_8__N_107[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_15.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_16 (.A(state[2]), .B(n42806), .C(n118[3]), 
         .Z(cur_pixel_8__N_107[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_16.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_17 (.A(state[2]), .B(n42806), .C(n118[2]), 
         .Z(cur_pixel_8__N_107[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_17.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_18 (.A(state[2]), .B(n42806), .C(n118[1]), 
         .Z(cur_pixel_8__N_107[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_18.init = 16'h1010;
    LUT4 i1_2_lut_rep_836 (.A(state[1]), .B(state[2]), .Z(n54839)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_836.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(n447[1]), 
         .D(state[0]), .Z(n71)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_rep_722_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n54725)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_rep_722_3_lut.init = 16'hefef;
    LUT4 i23033_4_lut (.A(sclk_c_enable_960), .B(n54725), .C(n6297), .D(n54609), 
         .Z(n35225)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i23033_4_lut.init = 16'haaa2;
    LUT4 i1_2_lut_3_lut_4_lut_adj_19 (.A(state[1]), .B(state[2]), .C(n447[0]), 
         .D(state[0]), .Z(n74)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_19.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_adj_20 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n14750[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_adj_20.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(n13381), 
         .Z(sclk_c_enable_71)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i1_3_lut_rep_735_4_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(sclk_c_enable_2472)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_3_lut_rep_735_4_lut_3_lut.init = 16'h8989;
    LUT4 i30309_2_lut_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .Z(n42478)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i30309_2_lut_3_lut.init = 16'hf8f8;
    LUT4 mux_1938_i1_4_lut (.A(n74), .B(n14750[0]), .C(n6297), .D(n52736), 
         .Z(n6298[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i1_4_lut.init = 16'hcfca;
    LUT4 i1950_3_lut (.A(state[2]), .B(state[1]), .C(n13381), .Z(n6297)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1950_3_lut.init = 16'ha8a8;
    LUT4 i8_4_lut (.A(n15), .B(cur_pixel[2]), .C(n14), .D(cur_pixel[3]), 
         .Z(n42806)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(cur_pixel[5]), .B(cur_pixel[1]), .C(cur_pixel[8]), 
         .D(cur_pixel[6]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i5_3_lut (.A(cur_pixel[4]), .B(cur_pixel[0]), .C(cur_pixel[7]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i5_3_lut.init = 16'h8080;
    LUT4 i38082_3_lut (.A(pixel[22]), .B(pixel[23]), .C(bit_counter[0]), 
         .Z(n53288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38082_3_lut.init = 16'hcaca;
    LUT4 i38081_3_lut (.A(pixel[20]), .B(pixel[21]), .C(bit_counter[0]), 
         .Z(n53287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38081_3_lut.init = 16'hcaca;
    LUT4 i38080_3_lut (.A(pixel[18]), .B(pixel[19]), .C(bit_counter[0]), 
         .Z(n53286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38080_3_lut.init = 16'hcaca;
    LUT4 i38079_3_lut (.A(pixel[16]), .B(pixel[17]), .C(bit_counter[0]), 
         .Z(n53285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38079_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut_adj_21 (.A(n54747), .B(state[1]), .C(n54663), 
         .D(n54664), .Z(n52736)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_3_lut_4_lut_4_lut_adj_21.init = 16'hce02;
    LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.A(state[0]), .B(n54839), .C(n13346), 
         .D(n42806), .Z(n9385[0])) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam i1_2_lut_3_lut_4_lut_adj_22.init = 16'hfddd;
    LUT4 mux_1928_i5_4_lut_4_lut (.A(state[0]), .B(n54839), .C(n447[4]), 
         .D(n54609), .Z(n6224[4])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !((D)+!C)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(42[12:17])
    defparam mux_1928_i5_4_lut_4_lut.init = 16'haad0;
    L6MUX21 i37834 (.D0(n53038), .D1(n53039), .SD(bit_counter[3]), .Z(n53040));
    PFUMX i38083 (.BLUT(n53285), .ALUT(n53286), .C0(bit_counter[1]), .Z(n53289));
    PFUMX i38084 (.BLUT(n53287), .ALUT(n53288), .C0(bit_counter[1]), .Z(n53290));
    LUT4 i37827_3_lut (.A(pixel[14]), .B(pixel[15]), .C(bit_counter[0]), 
         .Z(n53033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37827_3_lut.init = 16'hcaca;
    LUT4 i37826_3_lut (.A(pixel[12]), .B(pixel[13]), .C(bit_counter[0]), 
         .Z(n53032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37826_3_lut.init = 16'hcaca;
    LUT4 i37825_3_lut (.A(pixel[10]), .B(pixel[11]), .C(bit_counter[0]), 
         .Z(n53031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37825_3_lut.init = 16'hcaca;
    LUT4 i37824_3_lut (.A(pixel[8]), .B(pixel[9]), .C(bit_counter[0]), 
         .Z(n53030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37824_3_lut.init = 16'hcaca;
    LUT4 i37823_3_lut (.A(pixel[6]), .B(pixel[7]), .C(bit_counter[0]), 
         .Z(n53029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37823_3_lut.init = 16'hcaca;
    LUT4 i37822_3_lut (.A(pixel[4]), .B(pixel[5]), .C(bit_counter[0]), 
         .Z(n53028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37822_3_lut.init = 16'hcaca;
    LUT4 i37821_3_lut (.A(pixel[2]), .B(pixel[3]), .C(bit_counter[0]), 
         .Z(n53027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37821_3_lut.init = 16'hcaca;
    LUT4 i37820_3_lut (.A(pixel[0]), .B(pixel[1]), .C(bit_counter[0]), 
         .Z(n53026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37820_3_lut.init = 16'hcaca;
    CCU2D add_33922_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49102), 
          .S0(n13381));
    defparam add_33922_cout.INIT0 = 16'h0000;
    defparam add_33922_cout.INIT1 = 16'h0000;
    defparam add_33922_cout.INJECT1_0 = "NO";
    defparam add_33922_cout.INJECT1_1 = "NO";
    CCU2D add_33922_31 (.A0(delay_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49101), .COUT(n49102));
    defparam add_33922_31.INIT0 = 16'hf555;
    defparam add_33922_31.INIT1 = 16'h5555;
    defparam add_33922_31.INJECT1_0 = "NO";
    defparam add_33922_31.INJECT1_1 = "NO";
    CCU2D add_33922_29 (.A0(delay_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49100), .COUT(n49101));
    defparam add_33922_29.INIT0 = 16'hf555;
    defparam add_33922_29.INIT1 = 16'hf555;
    defparam add_33922_29.INJECT1_0 = "NO";
    defparam add_33922_29.INJECT1_1 = "NO";
    CCU2D add_33922_27 (.A0(delay_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49099), .COUT(n49100));
    defparam add_33922_27.INIT0 = 16'hf555;
    defparam add_33922_27.INIT1 = 16'hf555;
    defparam add_33922_27.INJECT1_0 = "NO";
    defparam add_33922_27.INJECT1_1 = "NO";
    CCU2D add_33922_25 (.A0(delay_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49098), .COUT(n49099));
    defparam add_33922_25.INIT0 = 16'hf555;
    defparam add_33922_25.INIT1 = 16'hf555;
    defparam add_33922_25.INJECT1_0 = "NO";
    defparam add_33922_25.INJECT1_1 = "NO";
    CCU2D add_33922_23 (.A0(delay_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49097), .COUT(n49098));
    defparam add_33922_23.INIT0 = 16'hf555;
    defparam add_33922_23.INIT1 = 16'hf555;
    defparam add_33922_23.INJECT1_0 = "NO";
    defparam add_33922_23.INJECT1_1 = "NO";
    CCU2D add_33922_21 (.A0(delay_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49096), .COUT(n49097));
    defparam add_33922_21.INIT0 = 16'hf555;
    defparam add_33922_21.INIT1 = 16'hf555;
    defparam add_33922_21.INJECT1_0 = "NO";
    defparam add_33922_21.INJECT1_1 = "NO";
    CCU2D add_33922_19 (.A0(delay_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49095), .COUT(n49096));
    defparam add_33922_19.INIT0 = 16'hf555;
    defparam add_33922_19.INIT1 = 16'hf555;
    defparam add_33922_19.INJECT1_0 = "NO";
    defparam add_33922_19.INJECT1_1 = "NO";
    CCU2D add_33922_17 (.A0(delay_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49094), .COUT(n49095));
    defparam add_33922_17.INIT0 = 16'hf555;
    defparam add_33922_17.INIT1 = 16'hf555;
    defparam add_33922_17.INJECT1_0 = "NO";
    defparam add_33922_17.INJECT1_1 = "NO";
    CCU2D add_33922_15 (.A0(delay_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49093), .COUT(n49094));
    defparam add_33922_15.INIT0 = 16'hf555;
    defparam add_33922_15.INIT1 = 16'hf555;
    defparam add_33922_15.INJECT1_0 = "NO";
    defparam add_33922_15.INJECT1_1 = "NO";
    CCU2D add_33922_13 (.A0(delay_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49092), .COUT(n49093));
    defparam add_33922_13.INIT0 = 16'hf555;
    defparam add_33922_13.INIT1 = 16'hf555;
    defparam add_33922_13.INJECT1_0 = "NO";
    defparam add_33922_13.INJECT1_1 = "NO";
    CCU2D add_33922_11 (.A0(delay_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49091), .COUT(n49092));
    defparam add_33922_11.INIT0 = 16'hf555;
    defparam add_33922_11.INIT1 = 16'hf555;
    defparam add_33922_11.INJECT1_0 = "NO";
    defparam add_33922_11.INJECT1_1 = "NO";
    CCU2D add_33922_9 (.A0(delay_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49090), .COUT(n49091));
    defparam add_33922_9.INIT0 = 16'hf555;
    defparam add_33922_9.INIT1 = 16'hf555;
    defparam add_33922_9.INJECT1_0 = "NO";
    defparam add_33922_9.INJECT1_1 = "NO";
    CCU2D add_33922_7 (.A0(delay_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49089), .COUT(n49090));
    defparam add_33922_7.INIT0 = 16'hf555;
    defparam add_33922_7.INIT1 = 16'hf555;
    defparam add_33922_7.INJECT1_0 = "NO";
    defparam add_33922_7.INJECT1_1 = "NO";
    CCU2D add_33922_5 (.A0(delay_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49088), .COUT(n49089));
    defparam add_33922_5.INIT0 = 16'hf555;
    defparam add_33922_5.INIT1 = 16'hf555;
    defparam add_33922_5.INJECT1_0 = "NO";
    defparam add_33922_5.INJECT1_1 = "NO";
    CCU2D add_33922_3 (.A0(delay_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49087), .COUT(n49088));
    defparam add_33922_3.INIT0 = 16'hf555;
    defparam add_33922_3.INIT1 = 16'hf555;
    defparam add_33922_3.INJECT1_0 = "NO";
    defparam add_33922_3.INJECT1_1 = "NO";
    CCU2D add_33922_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(delay_counter[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n49087));
    defparam add_33922_1.INIT0 = 16'hF000;
    defparam add_33922_1.INIT1 = 16'ha666;
    defparam add_33922_1.INJECT1_0 = "NO";
    defparam add_33922_1.INJECT1_1 = "NO";
    CCU2D add_33923_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n49086), 
          .S0(n13346));
    defparam add_33923_cout.INIT0 = 16'h0000;
    defparam add_33923_cout.INIT1 = 16'h0000;
    defparam add_33923_cout.INJECT1_0 = "NO";
    defparam add_33923_cout.INJECT1_1 = "NO";
    CCU2D add_33923_31 (.A0(bit_counter[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[31]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49085), .COUT(n49086));
    defparam add_33923_31.INIT0 = 16'hf555;
    defparam add_33923_31.INIT1 = 16'h5555;
    defparam add_33923_31.INJECT1_0 = "NO";
    defparam add_33923_31.INJECT1_1 = "NO";
    CCU2D add_33923_29 (.A0(bit_counter[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[29]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49084), .COUT(n49085));
    defparam add_33923_29.INIT0 = 16'hf555;
    defparam add_33923_29.INIT1 = 16'hf555;
    defparam add_33923_29.INJECT1_0 = "NO";
    defparam add_33923_29.INJECT1_1 = "NO";
    CCU2D add_33923_27 (.A0(bit_counter[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[27]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49083), .COUT(n49084));
    defparam add_33923_27.INIT0 = 16'hf555;
    defparam add_33923_27.INIT1 = 16'hf555;
    defparam add_33923_27.INJECT1_0 = "NO";
    defparam add_33923_27.INJECT1_1 = "NO";
    CCU2D add_33923_25 (.A0(bit_counter[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49082), .COUT(n49083));
    defparam add_33923_25.INIT0 = 16'hf555;
    defparam add_33923_25.INIT1 = 16'hf555;
    defparam add_33923_25.INJECT1_0 = "NO";
    defparam add_33923_25.INJECT1_1 = "NO";
    CCU2D add_33923_23 (.A0(bit_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49081), .COUT(n49082));
    defparam add_33923_23.INIT0 = 16'hf555;
    defparam add_33923_23.INIT1 = 16'hf555;
    defparam add_33923_23.INJECT1_0 = "NO";
    defparam add_33923_23.INJECT1_1 = "NO";
    CCU2D add_33923_21 (.A0(bit_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49080), .COUT(n49081));
    defparam add_33923_21.INIT0 = 16'hf555;
    defparam add_33923_21.INIT1 = 16'hf555;
    defparam add_33923_21.INJECT1_0 = "NO";
    defparam add_33923_21.INJECT1_1 = "NO";
    CCU2D add_33923_19 (.A0(bit_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49079), .COUT(n49080));
    defparam add_33923_19.INIT0 = 16'hf555;
    defparam add_33923_19.INIT1 = 16'hf555;
    defparam add_33923_19.INJECT1_0 = "NO";
    defparam add_33923_19.INJECT1_1 = "NO";
    CCU2D add_33923_17 (.A0(bit_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49078), .COUT(n49079));
    defparam add_33923_17.INIT0 = 16'hf555;
    defparam add_33923_17.INIT1 = 16'hf555;
    defparam add_33923_17.INJECT1_0 = "NO";
    defparam add_33923_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_744 (.A(state[2]), .B(state[0]), .Z(n54747)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_rep_744.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(state[2]), .B(state[0]), .C(n13346), 
         .D(state[1]), .Z(n39073)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h0004;
    LUT4 i11_3_lut (.A(state[0]), .B(state[2]), .C(state[1]), .Z(sclk_c_enable_70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    CCU2D add_33923_15 (.A0(bit_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49077), .COUT(n49078));
    defparam add_33923_15.INIT0 = 16'hf555;
    defparam add_33923_15.INIT1 = 16'hf555;
    defparam add_33923_15.INJECT1_0 = "NO";
    defparam add_33923_15.INJECT1_1 = "NO";
    LUT4 bit_counter_4__I_0_i31_4_lut (.A(n53040), .B(n53291), .C(bit_counter[4]), 
         .D(bit_counter[3]), .Z(serial_N_437)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(88[22:33])
    defparam bit_counter_4__I_0_i31_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_3_lut_adj_24 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[31]), 
         .Z(bit_counter_31__N_172[31])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_24.init = 16'h4040;
    CCU2D add_33923_13 (.A0(bit_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49076), .COUT(n49077));
    defparam add_33923_13.INIT0 = 16'hf555;
    defparam add_33923_13.INIT1 = 16'hf555;
    defparam add_33923_13.INJECT1_0 = "NO";
    defparam add_33923_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_25 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[30]), 
         .Z(bit_counter_31__N_172[30])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_25.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_26 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[29]), 
         .Z(bit_counter_31__N_172[29])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_26.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_27 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[28]), 
         .Z(bit_counter_31__N_172[28])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_27.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_28 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[27]), 
         .Z(bit_counter_31__N_172[27])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_28.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_29 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[26]), 
         .Z(bit_counter_31__N_172[26])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_29.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_30 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[25]), 
         .Z(bit_counter_31__N_172[25])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_30.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_31 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[24]), 
         .Z(bit_counter_31__N_172[24])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_31.init = 16'h4040;
    CCU2D add_33923_11 (.A0(bit_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49075), .COUT(n49076));
    defparam add_33923_11.INIT0 = 16'hf555;
    defparam add_33923_11.INIT1 = 16'hf555;
    defparam add_33923_11.INJECT1_0 = "NO";
    defparam add_33923_11.INJECT1_1 = "NO";
    LUT4 i29470_4_lut (.A(n9385[0]), .B(n9392), .C(state[0]), .D(n54651), 
         .Z(state_2__N_104[0])) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i29470_4_lut.init = 16'h0322;
    LUT4 i1_4_lut (.A(state[2]), .B(state[0]), .C(state[1]), .D(n13381), 
         .Z(n9392)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam i1_4_lut.init = 16'ha8a0;
    LUT4 i1_2_lut_3_lut_adj_32 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[23]), 
         .Z(bit_counter_31__N_172[23])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_32.init = 16'h4040;
    CCU2D add_33923_9 (.A0(bit_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49074), .COUT(n49075));
    defparam add_33923_9.INIT0 = 16'hf555;
    defparam add_33923_9.INIT1 = 16'hf555;
    defparam add_33923_9.INJECT1_0 = "NO";
    defparam add_33923_9.INJECT1_1 = "NO";
    CCU2D add_33923_7 (.A0(bit_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49073), .COUT(n49074));
    defparam add_33923_7.INIT0 = 16'hf555;
    defparam add_33923_7.INIT1 = 16'hf555;
    defparam add_33923_7.INJECT1_0 = "NO";
    defparam add_33923_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_33 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[22]), 
         .Z(bit_counter_31__N_172[22])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_33.init = 16'h4040;
    CCU2D add_33923_5 (.A0(bit_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49072), .COUT(n49073));
    defparam add_33923_5.INIT0 = 16'hf555;
    defparam add_33923_5.INIT1 = 16'hf555;
    defparam add_33923_5.INJECT1_0 = "NO";
    defparam add_33923_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_34 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[21]), 
         .Z(bit_counter_31__N_172[21])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_34.init = 16'h4040;
    CCU2D add_33923_3 (.A0(bit_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(bit_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n49071), .COUT(n49072));
    defparam add_33923_3.INIT0 = 16'hf555;
    defparam add_33923_3.INIT1 = 16'hf555;
    defparam add_33923_3.INJECT1_0 = "NO";
    defparam add_33923_3.INJECT1_1 = "NO";
    CCU2D add_33923_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(bit_counter[0]), .B1(bit_counter[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n49071));
    defparam add_33923_1.INIT0 = 16'hF000;
    defparam add_33923_1.INIT1 = 16'ha666;
    defparam add_33923_1.INJECT1_0 = "NO";
    defparam add_33923_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_35 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[20]), 
         .Z(bit_counter_31__N_172[20])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_35.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_36 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[19]), 
         .Z(bit_counter_31__N_172[19])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_36.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_37 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[18]), 
         .Z(bit_counter_31__N_172[18])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_37.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_38 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[17]), 
         .Z(bit_counter_31__N_172[17])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_38.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_39 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[16]), 
         .Z(bit_counter_31__N_172[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_39.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_40 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[15]), 
         .Z(bit_counter_31__N_172[15])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_40.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_41 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[14]), 
         .Z(bit_counter_31__N_172[14])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_41.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_42 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[13]), 
         .Z(bit_counter_31__N_172[13])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_42.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_43 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[12]), 
         .Z(bit_counter_31__N_172[12])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_43.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_44 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[11]), 
         .Z(bit_counter_31__N_172[11])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_44.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_45 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[10]), 
         .Z(bit_counter_31__N_172[10])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_45.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_46 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[9]), 
         .Z(bit_counter_31__N_172[9])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_46.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_47 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[8]), 
         .Z(bit_counter_31__N_172[8])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_47.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_48 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[7]), 
         .Z(bit_counter_31__N_172[7])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_48.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_49 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[6]), 
         .Z(bit_counter_31__N_172[6])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_49.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_50 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[5]), 
         .Z(bit_counter_31__N_172[5])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_50.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_51 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[2]), 
         .Z(bit_counter_31__N_172[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_51.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_52 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[1]), 
         .Z(bit_counter_31__N_172[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_52.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_53 (.A(state[2]), .B(state[0]), .C(bit_counter_31__N_204[0]), 
         .Z(bit_counter_31__N_172[0])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_2_lut_3_lut_adj_53.init = 16'h4040;
    LUT4 i38398_2_lut_rep_745 (.A(state[2]), .B(state[1]), .Z(sclk_c_enable_1182)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i38398_2_lut_rep_745.init = 16'h9999;
    LUT4 i23162_2_lut_2_lut (.A(state[2]), .B(state[1]), .Z(n35403)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23162_2_lut_2_lut.init = 16'h8888;
    CCU2D add_50_33 (.A0(delay_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47729), .S0(n447[31]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_33.INIT0 = 16'h5555;
    defparam add_50_33.INIT1 = 16'h0000;
    defparam add_50_33.INJECT1_0 = "NO";
    defparam add_50_33.INJECT1_1 = "NO";
    CCU2D add_50_31 (.A0(delay_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47728), .COUT(n47729), .S0(n447[29]), 
          .S1(n447[30]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_31.INIT0 = 16'h5555;
    defparam add_50_31.INIT1 = 16'h5555;
    defparam add_50_31.INJECT1_0 = "NO";
    defparam add_50_31.INJECT1_1 = "NO";
    CCU2D add_50_29 (.A0(delay_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47727), .COUT(n47728), .S0(n447[27]), 
          .S1(n447[28]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_29.INIT0 = 16'h5555;
    defparam add_50_29.INIT1 = 16'h5555;
    defparam add_50_29.INJECT1_0 = "NO";
    defparam add_50_29.INJECT1_1 = "NO";
    LUT4 i28770_2_lut (.A(bit_counter_31__N_204[4]), .B(state[0]), .Z(n1)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28770_2_lut.init = 16'hbbbb;
    CCU2D add_50_27 (.A0(delay_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47726), .COUT(n47727), .S0(n447[25]), 
          .S1(n447[26]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_27.INIT0 = 16'h5555;
    defparam add_50_27.INIT1 = 16'h5555;
    defparam add_50_27.INJECT1_0 = "NO";
    defparam add_50_27.INJECT1_1 = "NO";
    LUT4 i28769_2_lut (.A(bit_counter_31__N_204[3]), .B(state[0]), .Z(n1_adj_895)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i28769_2_lut.init = 16'hbbbb;
    CCU2D add_50_25 (.A0(delay_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47725), .COUT(n47726), .S0(n447[23]), 
          .S1(n447[24]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_25.INIT0 = 16'h5555;
    defparam add_50_25.INIT1 = 16'h5555;
    defparam add_50_25.INJECT1_0 = "NO";
    defparam add_50_25.INJECT1_1 = "NO";
    CCU2D add_50_23 (.A0(delay_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47724), .COUT(n47725), .S0(n447[21]), 
          .S1(n447[22]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_23.INIT0 = 16'h5555;
    defparam add_50_23.INIT1 = 16'h5555;
    defparam add_50_23.INJECT1_0 = "NO";
    defparam add_50_23.INJECT1_1 = "NO";
    CCU2D add_50_21 (.A0(delay_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47723), .COUT(n47724), .S0(n447[19]), 
          .S1(n447[20]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_21.INIT0 = 16'h5555;
    defparam add_50_21.INIT1 = 16'h5555;
    defparam add_50_21.INJECT1_0 = "NO";
    defparam add_50_21.INJECT1_1 = "NO";
    CCU2D add_50_19 (.A0(delay_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47722), .COUT(n47723), .S0(n447[17]), 
          .S1(n447[18]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_19.INIT0 = 16'h5555;
    defparam add_50_19.INIT1 = 16'h5555;
    defparam add_50_19.INJECT1_0 = "NO";
    defparam add_50_19.INJECT1_1 = "NO";
    CCU2D add_50_17 (.A0(delay_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47721), .COUT(n47722), .S0(n447[15]), 
          .S1(n447[16]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_17.INIT0 = 16'h5555;
    defparam add_50_17.INIT1 = 16'h5555;
    defparam add_50_17.INJECT1_0 = "NO";
    defparam add_50_17.INJECT1_1 = "NO";
    CCU2D add_50_15 (.A0(delay_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47720), .COUT(n47721), .S0(n447[13]), 
          .S1(n447[14]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_15.INIT0 = 16'h5555;
    defparam add_50_15.INIT1 = 16'h5555;
    defparam add_50_15.INJECT1_0 = "NO";
    defparam add_50_15.INJECT1_1 = "NO";
    CCU2D add_50_13 (.A0(delay_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47719), .COUT(n47720), .S0(n447[11]), 
          .S1(n447[12]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_13.INIT0 = 16'h5555;
    defparam add_50_13.INIT1 = 16'h5555;
    defparam add_50_13.INJECT1_0 = "NO";
    defparam add_50_13.INJECT1_1 = "NO";
    CCU2D add_50_11 (.A0(delay_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47718), .COUT(n47719), .S0(n447[9]), .S1(n447[10]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_11.INIT0 = 16'h5555;
    defparam add_50_11.INIT1 = 16'h5555;
    defparam add_50_11.INJECT1_0 = "NO";
    defparam add_50_11.INJECT1_1 = "NO";
    CCU2D add_50_9 (.A0(delay_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47717), .COUT(n47718), .S0(n447[7]), .S1(n447[8]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_9.INIT0 = 16'h5555;
    defparam add_50_9.INIT1 = 16'h5555;
    defparam add_50_9.INJECT1_0 = "NO";
    defparam add_50_9.INJECT1_1 = "NO";
    CCU2D add_50_7 (.A0(delay_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47716), .COUT(n47717), .S0(n447[5]), .S1(n447[6]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_7.INIT0 = 16'h5555;
    defparam add_50_7.INIT1 = 16'h5555;
    defparam add_50_7.INJECT1_0 = "NO";
    defparam add_50_7.INJECT1_1 = "NO";
    CCU2D add_50_5 (.A0(delay_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47715), .COUT(n47716), .S0(n447[3]), .S1(n447[4]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_5.INIT0 = 16'h5555;
    defparam add_50_5.INIT1 = 16'h5555;
    defparam add_50_5.INJECT1_0 = "NO";
    defparam add_50_5.INJECT1_1 = "NO";
    CCU2D add_50_3 (.A0(delay_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n47714), .COUT(n47715), .S0(n447[1]), .S1(n447[2]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_3.INIT0 = 16'h5555;
    defparam add_50_3.INIT1 = 16'h5555;
    defparam add_50_3.INJECT1_0 = "NO";
    defparam add_50_3.INJECT1_1 = "NO";
    LUT4 i23009_2_lut_4_lut (.A(n54664), .B(state[0]), .C(state[1]), .D(n6297), 
         .Z(n35221)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i23009_2_lut_4_lut.init = 16'hfd00;
    CCU2D add_50_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47714), .S1(n447[0]));   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(106[23:36])
    defparam add_50_1.INIT0 = 16'hF000;
    defparam add_50_1.INIT1 = 16'h5555;
    defparam add_50_1.INJECT1_0 = "NO";
    defparam add_50_1.INJECT1_1 = "NO";
    CCU2D add_17_9 (.A0(cur_pixel[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47712), .S0(n118[7]), .S1(n118[8]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_9.INIT0 = 16'h5aaa;
    defparam add_17_9.INIT1 = 16'h5aaa;
    defparam add_17_9.INJECT1_0 = "NO";
    defparam add_17_9.INJECT1_1 = "NO";
    CCU2D add_17_7 (.A0(cur_pixel[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47711), .COUT(n47712), .S0(n118[5]), .S1(n118[6]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_7.INIT0 = 16'h5aaa;
    defparam add_17_7.INIT1 = 16'h5aaa;
    defparam add_17_7.INJECT1_0 = "NO";
    defparam add_17_7.INJECT1_1 = "NO";
    LUT4 mux_1938_i2_4_lut (.A(n71), .B(n14750[0]), .C(n6297), .D(n52736), 
         .Z(n6298[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i2_4_lut.init = 16'hcfca;
    LUT4 mux_1938_i4_4_lut (.A(n39073), .B(n42478), .C(n6297), .D(n4), 
         .Z(n6298[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i4_4_lut.init = 16'h3f3a;
    LUT4 i1_4_lut_adj_54 (.A(n42806), .B(n54609), .C(n447[3]), .D(n54725), 
         .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam i1_4_lut_adj_54.init = 16'hfcee;
    CCU2D add_17_5 (.A0(cur_pixel[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47710), .COUT(n47711), .S0(n118[3]), .S1(n118[4]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_5.INIT0 = 16'h5aaa;
    defparam add_17_5.INIT1 = 16'h5aaa;
    defparam add_17_5.INJECT1_0 = "NO";
    defparam add_17_5.INJECT1_1 = "NO";
    LUT4 mux_1938_i8_4_lut (.A(n6122[7]), .B(n42478), .C(n6297), .D(n54609), 
         .Z(n6298[7])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i8_4_lut.init = 16'h303a;
    FD1P3IX pixel_i23 (.D(\Q[7] [23]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i23.GSR = "DISABLED";
    FD1P3IX pixel_i22 (.D(\Q[7] [22]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i22.GSR = "DISABLED";
    CCU2D add_17_3 (.A0(cur_pixel[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n47709), .COUT(n47710), .S0(n118[1]), .S1(n118[2]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_3.INIT0 = 16'h5aaa;
    defparam add_17_3.INIT1 = 16'h5aaa;
    defparam add_17_3.INJECT1_0 = "NO";
    defparam add_17_3.INJECT1_1 = "NO";
    FD1P3IX pixel_i21 (.D(\Q[7] [21]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i21.GSR = "DISABLED";
    FD1P3IX pixel_i20 (.D(\Q[7] [20]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i20.GSR = "DISABLED";
    FD1P3IX pixel_i19 (.D(\Q[7] [19]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i19.GSR = "DISABLED";
    FD1P3IX pixel_i18 (.D(\Q[7] [18]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i18.GSR = "DISABLED";
    LUT4 mux_1938_i9_4_lut (.A(n6122[8]), .B(n42478), .C(n6297), .D(n54609), 
         .Z(n6298[8])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i9_4_lut.init = 16'h303a;
    LUT4 mux_1938_i10_4_lut (.A(n80), .B(n42478), .C(n6297), .D(n54609), 
         .Z(n6298[9])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i10_4_lut.init = 16'h303a;
    CCU2D add_17_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cur_pixel[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n47709), .S1(n118[0]));   // C:/lscc/diamond/3.13/ispfpga/vhdl_packages/syn_unsi.vhd(118[20:31])
    defparam add_17_1.INIT0 = 16'hF000;
    defparam add_17_1.INIT1 = 16'h5555;
    defparam add_17_1.INJECT1_0 = "NO";
    defparam add_17_1.INJECT1_1 = "NO";
    LUT4 mux_1938_i13_4_lut (.A(n6122[12]), .B(n42478), .C(n6297), .D(n54609), 
         .Z(n6298[12])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(51[3] 113[12])
    defparam mux_1938_i13_4_lut.init = 16'h303a;
    FD1P3IX pixel_i17 (.D(\Q[7] [17]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i17.GSR = "DISABLED";
    FD1P3IX pixel_i16 (.D(\Q[7] [16]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i16.GSR = "DISABLED";
    FD1P3IX pixel_i15 (.D(\Q[7] [15]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i15.GSR = "DISABLED";
    FD1P3IX pixel_i14 (.D(\Q[7] [14]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i14.GSR = "DISABLED";
    FD1P3IX pixel_i13 (.D(\Q[7] [13]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i13.GSR = "DISABLED";
    FD1P3IX pixel_i12 (.D(\Q[7] [12]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i12.GSR = "DISABLED";
    FD1P3IX pixel_i11 (.D(\Q[7] [11]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i11.GSR = "DISABLED";
    FD1P3IX pixel_i10 (.D(\Q[7] [10]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i10.GSR = "DISABLED";
    FD1P3IX pixel_i9 (.D(\Q[7] [9]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i9.GSR = "DISABLED";
    FD1P3IX pixel_i8 (.D(\Q[7] [8]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i8.GSR = "DISABLED";
    FD1P3IX pixel_i7 (.D(\Q[7] [7]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i7.GSR = "DISABLED";
    FD1P3IX pixel_i6 (.D(\Q[7] [6]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i6.GSR = "DISABLED";
    FD1P3IX pixel_i5 (.D(\Q[7] [5]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i5.GSR = "DISABLED";
    FD1P3IX pixel_i4 (.D(\Q[7] [4]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i4.GSR = "DISABLED";
    FD1P3IX pixel_i3 (.D(\Q[7] [3]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i3.GSR = "DISABLED";
    FD1P3IX pixel_i2 (.D(\Q[7] [2]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i2.GSR = "DISABLED";
    FD1P3IX pixel_i1 (.D(\Q[7] [1]), .SP(sclk_c_enable_2472), .CD(n35403), 
            .CK(sclk_c), .Q(pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam pixel_i1.GSR = "DISABLED";
    FD1P3AX cur_pixel_i8 (.D(cur_pixel_8__N_107[8]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i8.GSR = "DISABLED";
    FD1P3AX cur_pixel_i7 (.D(cur_pixel_8__N_107[7]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i7.GSR = "DISABLED";
    FD1P3AX cur_pixel_i6 (.D(cur_pixel_8__N_107[6]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i6.GSR = "DISABLED";
    FD1P3AX cur_pixel_i5 (.D(cur_pixel_8__N_107[5]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i5.GSR = "DISABLED";
    FD1P3AX cur_pixel_i4 (.D(cur_pixel_8__N_107[4]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i4.GSR = "DISABLED";
    FD1P3AX cur_pixel_i3 (.D(cur_pixel_8__N_107[3]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i3.GSR = "DISABLED";
    FD1P3AX cur_pixel_i2 (.D(cur_pixel_8__N_107[2]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i2.GSR = "DISABLED";
    FD1P3AX cur_pixel_i1 (.D(cur_pixel_8__N_107[1]), .SP(sclk_c_enable_2480), 
            .CK(sclk_c), .Q(cur_pixel[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=12, LSE_RCOL=18, LSE_LLINE=212, LSE_RLINE=212 */ ;   // c:/users/ryanm/onedrive/documents/diamond/ws2812_driver/xo3d/source/ws2812.vhd(41[2] 114[14])
    defparam cur_pixel_i1.GSR = "DISABLED";
    PFUMX i38963 (.BLUT(n54983), .ALUT(n54984), .C0(state[1]), .Z(n54985));
    PFUMX i38913 (.BLUT(n54907), .ALUT(n54908), .C0(state[1]), .Z(state_2__N_104[1]));
    
endmodule
